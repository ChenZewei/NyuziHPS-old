// fpga_sdram_controller.v

// Generated using ACDS version 13.0sp1 232 at 2015.08.06.11:37:57

`timescale 1 ps / 1 ps
module fpga_sdram_controller (
		input  wire        clk_clk,              //      clk.clk
		input  wire        reset_reset_n,        //    reset.reset_n
		output wire [12:0] memory_mem_a,         //   memory.mem_a
		output wire [2:0]  memory_mem_ba,        //         .mem_ba
		output wire [0:0]  memory_mem_ck,        //         .mem_ck
		output wire [0:0]  memory_mem_ck_n,      //         .mem_ck_n
		output wire [0:0]  memory_mem_cke,       //         .mem_cke
		output wire [0:0]  memory_mem_cs_n,      //         .mem_cs_n
		output wire [0:0]  memory_mem_dm,        //         .mem_dm
		output wire [0:0]  memory_mem_ras_n,     //         .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,     //         .mem_cas_n
		output wire [0:0]  memory_mem_we_n,      //         .mem_we_n
		output wire        memory_mem_reset_n,   //         .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,        //         .mem_dq
		inout  wire [0:0]  memory_mem_dqs,       //         .mem_dqs
		inout  wire [0:0]  memory_mem_dqs_n,     //         .mem_dqs_n
		output wire [0:0]  memory_mem_odt,       //         .mem_odt
		input  wire        oct_rzqin,            //      oct.rzqin
		output wire [12:0] memory_0_mem_a,       // memory_0.mem_a
		output wire [2:0]  memory_0_mem_ba,      //         .mem_ba
		output wire        memory_0_mem_ck,      //         .mem_ck
		output wire        memory_0_mem_ck_n,    //         .mem_ck_n
		output wire        memory_0_mem_cke,     //         .mem_cke
		output wire        memory_0_mem_cs_n,    //         .mem_cs_n
		output wire        memory_0_mem_ras_n,   //         .mem_ras_n
		output wire        memory_0_mem_cas_n,   //         .mem_cas_n
		output wire        memory_0_mem_we_n,    //         .mem_we_n
		output wire        memory_0_mem_reset_n, //         .mem_reset_n
		inout  wire [7:0]  memory_0_mem_dq,      //         .mem_dq
		inout  wire        memory_0_mem_dqs,     //         .mem_dqs
		inout  wire        memory_0_mem_dqs_n,   //         .mem_dqs_n
		output wire        memory_0_mem_odt,     //         .mem_odt
		output wire        memory_0_mem_dm,      //         .mem_dm
		input  wire        memory_0_oct_rzqin    //         .oct_rzqin
	);

	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest;                           // mem_if_ddr3_emif_0:avl_ready -> mem_if_ddr3_emif_0_avl_translator:av_waitrequest
	wire    [5:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount;                            // mem_if_ddr3_emif_0_avl_translator:av_burstcount -> mem_if_ddr3_emif_0:avl_size
	wire   [31:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata;                             // mem_if_ddr3_emif_0_avl_translator:av_writedata -> mem_if_ddr3_emif_0:avl_wdata
	wire   [20:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address;                               // mem_if_ddr3_emif_0_avl_translator:av_address -> mem_if_ddr3_emif_0:avl_addr
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write;                                 // mem_if_ddr3_emif_0_avl_translator:av_write -> mem_if_ddr3_emif_0:avl_write_req
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer;                    // mem_if_ddr3_emif_0_avl_translator:av_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read;                                  // mem_if_ddr3_emif_0_avl_translator:av_read -> mem_if_ddr3_emif_0:avl_read_req
	wire   [31:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata;                              // mem_if_ddr3_emif_0:avl_rdata -> mem_if_ddr3_emif_0_avl_translator:av_readdata
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid;                         // mem_if_ddr3_emif_0:avl_rdata_valid -> mem_if_ddr3_emif_0_avl_translator:av_readdatavalid
	wire    [3:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable;                            // mem_if_ddr3_emif_0_avl_translator:av_byteenable -> mem_if_ddr3_emif_0:avl_be
	wire          mem_if_ddr3_emif_0_afi_clk_clk;                                                              // mem_if_ddr3_emif_0:afi_clk -> [burst_adapter:clk, cmd_xbar_mux:clk, crosser:out_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, id_router:clk, mem_if_ddr3_emif_0_avl_translator:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rst_controller:clk, width_adapter:clk]
	wire          hps_0_h2f_axi_master_awvalid;                                                                // hps_0:h2f_AWVALID -> hps_0_h2f_axi_master_agent:awvalid
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                                                 // hps_0:h2f_ARSIZE -> hps_0_h2f_axi_master_agent:arsize
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                                                 // hps_0:h2f_ARLOCK -> hps_0_h2f_axi_master_agent:arlock
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                                                // hps_0:h2f_AWCACHE -> hps_0_h2f_axi_master_agent:awcache
	wire          hps_0_h2f_axi_master_arready;                                                                // hps_0_h2f_axi_master_agent:arready -> hps_0:h2f_ARREADY
	wire   [11:0] hps_0_h2f_axi_master_arid;                                                                   // hps_0:h2f_ARID -> hps_0_h2f_axi_master_agent:arid
	wire          hps_0_h2f_axi_master_rready;                                                                 // hps_0:h2f_RREADY -> hps_0_h2f_axi_master_agent:rready
	wire          hps_0_h2f_axi_master_bready;                                                                 // hps_0:h2f_BREADY -> hps_0_h2f_axi_master_agent:bready
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                                                 // hps_0:h2f_AWSIZE -> hps_0_h2f_axi_master_agent:awsize
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                                                 // hps_0:h2f_AWPROT -> hps_0_h2f_axi_master_agent:awprot
	wire          hps_0_h2f_axi_master_arvalid;                                                                // hps_0:h2f_ARVALID -> hps_0_h2f_axi_master_agent:arvalid
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                                                 // hps_0:h2f_ARPROT -> hps_0_h2f_axi_master_agent:arprot
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                                    // hps_0_h2f_axi_master_agent:bid -> hps_0:h2f_BID
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                                                  // hps_0:h2f_ARLEN -> hps_0_h2f_axi_master_agent:arlen
	wire          hps_0_h2f_axi_master_awready;                                                                // hps_0_h2f_axi_master_agent:awready -> hps_0:h2f_AWREADY
	wire   [11:0] hps_0_h2f_axi_master_awid;                                                                   // hps_0:h2f_AWID -> hps_0_h2f_axi_master_agent:awid
	wire          hps_0_h2f_axi_master_bvalid;                                                                 // hps_0_h2f_axi_master_agent:bvalid -> hps_0:h2f_BVALID
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                                    // hps_0:h2f_WID -> hps_0_h2f_axi_master_agent:wid
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                                                 // hps_0:h2f_AWLOCK -> hps_0_h2f_axi_master_agent:awlock
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                                                // hps_0:h2f_AWBURST -> hps_0_h2f_axi_master_agent:awburst
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                                                  // hps_0_h2f_axi_master_agent:bresp -> hps_0:h2f_BRESP
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                                                  // hps_0:h2f_WSTRB -> hps_0_h2f_axi_master_agent:wstrb
	wire          hps_0_h2f_axi_master_rvalid;                                                                 // hps_0_h2f_axi_master_agent:rvalid -> hps_0:h2f_RVALID
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                                                  // hps_0:h2f_WDATA -> hps_0_h2f_axi_master_agent:wdata
	wire          hps_0_h2f_axi_master_wready;                                                                 // hps_0_h2f_axi_master_agent:wready -> hps_0:h2f_WREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                                                // hps_0:h2f_ARBURST -> hps_0_h2f_axi_master_agent:arburst
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                                                  // hps_0_h2f_axi_master_agent:rdata -> hps_0:h2f_RDATA
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                                                 // hps_0:h2f_ARADDR -> hps_0_h2f_axi_master_agent:araddr
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                                                // hps_0:h2f_ARCACHE -> hps_0_h2f_axi_master_agent:arcache
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                                                  // hps_0:h2f_AWLEN -> hps_0_h2f_axi_master_agent:awlen
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                                                 // hps_0:h2f_AWADDR -> hps_0_h2f_axi_master_agent:awaddr
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                                    // hps_0_h2f_axi_master_agent:rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_wvalid;                                                                 // hps_0:h2f_WVALID -> hps_0_h2f_axi_master_agent:wvalid
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                                                  // hps_0_h2f_axi_master_agent:rresp -> hps_0:h2f_RRESP
	wire          hps_0_h2f_axi_master_wlast;                                                                  // hps_0:h2f_WLAST -> hps_0_h2f_axi_master_agent:wlast
	wire          hps_0_h2f_axi_master_rlast;                                                                  // hps_0_h2f_axi_master_agent:rlast -> hps_0:h2f_RLAST
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // mem_if_ddr3_emif_0_avl_translator:uav_waitrequest -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [7:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> mem_if_ddr3_emif_0_avl_translator:uav_burstcount
	wire   [31:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata;               // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> mem_if_ddr3_emif_0_avl_translator:uav_writedata
	wire   [29:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address;                 // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_address -> mem_if_ddr3_emif_0_avl_translator:uav_address
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write;                   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_write -> mem_if_ddr3_emif_0_avl_translator:uav_write
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_lock -> mem_if_ddr3_emif_0_avl_translator:uav_lock
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_read -> mem_if_ddr3_emif_0_avl_translator:uav_read
	wire   [31:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                // mem_if_ddr3_emif_0_avl_translator:uav_readdata -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // mem_if_ddr3_emif_0_avl_translator:uav_readdatavalid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mem_if_ddr3_emif_0_avl_translator:uav_debugaccess
	wire    [3:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> mem_if_ddr3_emif_0_avl_translator:uav_byteenable
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [120:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [120:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          hps_0_h2f_axi_master_agent_write_cp_endofpacket;                                             // hps_0_h2f_axi_master_agent:write_cp_endofpacket -> addr_router:sink_endofpacket
	wire          hps_0_h2f_axi_master_agent_write_cp_valid;                                                   // hps_0_h2f_axi_master_agent:write_cp_valid -> addr_router:sink_valid
	wire          hps_0_h2f_axi_master_agent_write_cp_startofpacket;                                           // hps_0_h2f_axi_master_agent:write_cp_startofpacket -> addr_router:sink_startofpacket
	wire  [155:0] hps_0_h2f_axi_master_agent_write_cp_data;                                                    // hps_0_h2f_axi_master_agent:write_cp_data -> addr_router:sink_data
	wire          hps_0_h2f_axi_master_agent_write_cp_ready;                                                   // addr_router:sink_ready -> hps_0_h2f_axi_master_agent:write_cp_ready
	wire          hps_0_h2f_axi_master_agent_read_cp_endofpacket;                                              // hps_0_h2f_axi_master_agent:read_cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          hps_0_h2f_axi_master_agent_read_cp_valid;                                                    // hps_0_h2f_axi_master_agent:read_cp_valid -> addr_router_001:sink_valid
	wire          hps_0_h2f_axi_master_agent_read_cp_startofpacket;                                            // hps_0_h2f_axi_master_agent:read_cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [155:0] hps_0_h2f_axi_master_agent_read_cp_data;                                                     // hps_0_h2f_axi_master_agent:read_cp_data -> addr_router_001:sink_data
	wire          hps_0_h2f_axi_master_agent_read_cp_ready;                                                    // addr_router_001:sink_ready -> hps_0_h2f_axi_master_agent:read_cp_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid;                   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [119:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                           // burst_adapter:source0_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                 // burst_adapter:source0_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                         // burst_adapter:source0_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [119:0] burst_adapter_source0_data;                                                                  // burst_adapter:source0_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                 // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                               // burst_adapter:source0_channel -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          width_adapter_cmd_source_endofpacket;                                                        // width_adapter:cmd_out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_cmd_source_valid;                                                              // width_adapter:cmd_out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_cmd_source_startofpacket;                                                      // width_adapter:cmd_out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [119:0] width_adapter_cmd_source_data;                                                               // width_adapter:cmd_out_data -> burst_adapter:sink0_data
	wire    [1:0] width_adapter_cmd_source_channel;                                                            // width_adapter:cmd_out_channel -> burst_adapter:sink0_channel
	wire          width_adapter_cmd_source_ready;                                                              // burst_adapter:sink0_ready -> width_adapter:cmd_out_ready
	wire          id_router_src_endofpacket;                                                                   // id_router:src_endofpacket -> width_adapter:rsp_in_endofpacket
	wire          id_router_src_valid;                                                                         // id_router:src_valid -> width_adapter:rsp_in_valid
	wire          id_router_src_startofpacket;                                                                 // id_router:src_startofpacket -> width_adapter:rsp_in_startofpacket
	wire  [119:0] id_router_src_data;                                                                          // id_router:src_data -> width_adapter:rsp_in_data
	wire    [1:0] id_router_src_channel;                                                                       // id_router:src_channel -> width_adapter:rsp_in_channel
	wire          id_router_src_ready;                                                                         // width_adapter:rsp_in_ready -> id_router:src_ready
	wire          rst_controller_reset_out_reset;                                                              // rst_controller:reset_out -> [burst_adapter:reset, cmd_xbar_mux:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, id_router:reset, mem_if_ddr3_emif_0_avl_translator:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, width_adapter:reset]
	wire          mem_if_ddr3_emif_0_afi_reset_reset;                                                          // mem_if_ddr3_emif_0:afi_reset_n -> rst_controller:reset_in0
	wire          rst_controller_001_reset_out_reset;                                                          // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, hps_0_h2f_axi_master_agent:aresetn]
	wire          hps_0_h2f_reset_reset;                                                                       // hps_0:h2f_rst_n -> rst_controller_001:reset_in0
	wire          addr_router_src_endofpacket;                                                                 // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                       // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                               // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [155:0] addr_router_src_data;                                                                        // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] addr_router_src_channel;                                                                     // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                       // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          crosser_002_out_ready;                                                                       // hps_0_h2f_axi_master_agent:write_rp_ready -> crosser_002:out_ready
	wire          addr_router_001_src_endofpacket;                                                             // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                   // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                           // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [155:0] addr_router_001_src_data;                                                                    // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [1:0] addr_router_001_src_channel;                                                                 // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                   // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          crosser_003_out_ready;                                                                       // hps_0_h2f_axi_master_agent:read_rp_ready -> crosser_003:out_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                // cmd_xbar_mux:src_endofpacket -> width_adapter:cmd_in_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                      // cmd_xbar_mux:src_valid -> width_adapter:cmd_in_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                              // cmd_xbar_mux:src_startofpacket -> width_adapter:cmd_in_startofpacket
	wire  [155:0] cmd_xbar_mux_src_data;                                                                       // cmd_xbar_mux:src_data -> width_adapter:cmd_in_data
	wire    [1:0] cmd_xbar_mux_src_channel;                                                                    // cmd_xbar_mux:src_channel -> width_adapter:cmd_in_channel
	wire          cmd_xbar_mux_src_ready;                                                                      // width_adapter:cmd_in_ready -> cmd_xbar_mux:src_ready
	wire          width_adapter_rsp_source_endofpacket;                                                        // width_adapter:rsp_out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_rsp_source_valid;                                                              // width_adapter:rsp_out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_rsp_source_startofpacket;                                                      // width_adapter:rsp_out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [155:0] width_adapter_rsp_source_data;                                                               // width_adapter:rsp_out_data -> rsp_xbar_demux:sink_data
	wire    [1:0] width_adapter_rsp_source_channel;                                                            // width_adapter:rsp_out_channel -> rsp_xbar_demux:sink_channel
	wire          width_adapter_rsp_source_ready;                                                              // rsp_xbar_demux:sink_ready -> width_adapter:rsp_out_ready
	wire          crosser_out_endofpacket;                                                                     // crosser:out_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          crosser_out_valid;                                                                           // crosser:out_valid -> cmd_xbar_mux:sink0_valid
	wire          crosser_out_startofpacket;                                                                   // crosser:out_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [155:0] crosser_out_data;                                                                            // crosser:out_data -> cmd_xbar_mux:sink0_data
	wire    [1:0] crosser_out_channel;                                                                         // crosser:out_channel -> cmd_xbar_mux:sink0_channel
	wire          crosser_out_ready;                                                                           // cmd_xbar_mux:sink0_ready -> crosser:out_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                             // cmd_xbar_demux:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                   // cmd_xbar_demux:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                           // cmd_xbar_demux:src0_startofpacket -> crosser:in_startofpacket
	wire  [155:0] cmd_xbar_demux_src0_data;                                                                    // cmd_xbar_demux:src0_data -> crosser:in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                                 // cmd_xbar_demux:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                                   // crosser:in_ready -> cmd_xbar_demux:src0_ready
	wire          crosser_001_out_endofpacket;                                                                 // crosser_001:out_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          crosser_001_out_valid;                                                                       // crosser_001:out_valid -> cmd_xbar_mux:sink1_valid
	wire          crosser_001_out_startofpacket;                                                               // crosser_001:out_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [155:0] crosser_001_out_data;                                                                        // crosser_001:out_data -> cmd_xbar_mux:sink1_data
	wire    [1:0] crosser_001_out_channel;                                                                     // crosser_001:out_channel -> cmd_xbar_mux:sink1_channel
	wire          crosser_001_out_ready;                                                                       // cmd_xbar_mux:sink1_ready -> crosser_001:out_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                         // cmd_xbar_demux_001:src0_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                               // cmd_xbar_demux_001:src0_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                       // cmd_xbar_demux_001:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [155:0] cmd_xbar_demux_001_src0_data;                                                                // cmd_xbar_demux_001:src0_data -> crosser_001:in_data
	wire    [1:0] cmd_xbar_demux_001_src0_channel;                                                             // cmd_xbar_demux_001:src0_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                               // crosser_001:in_ready -> cmd_xbar_demux_001:src0_ready
	wire          crosser_002_out_endofpacket;                                                                 // crosser_002:out_endofpacket -> hps_0_h2f_axi_master_agent:write_rp_endofpacket
	wire          crosser_002_out_valid;                                                                       // crosser_002:out_valid -> hps_0_h2f_axi_master_agent:write_rp_valid
	wire          crosser_002_out_startofpacket;                                                               // crosser_002:out_startofpacket -> hps_0_h2f_axi_master_agent:write_rp_startofpacket
	wire  [155:0] crosser_002_out_data;                                                                        // crosser_002:out_data -> hps_0_h2f_axi_master_agent:write_rp_data
	wire    [1:0] crosser_002_out_channel;                                                                     // crosser_002:out_channel -> hps_0_h2f_axi_master_agent:write_rp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                             // rsp_xbar_demux:src0_endofpacket -> crosser_002:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                   // rsp_xbar_demux:src0_valid -> crosser_002:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                           // rsp_xbar_demux:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [155:0] rsp_xbar_demux_src0_data;                                                                    // rsp_xbar_demux:src0_data -> crosser_002:in_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                                 // rsp_xbar_demux:src0_channel -> crosser_002:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                                   // crosser_002:in_ready -> rsp_xbar_demux:src0_ready
	wire          crosser_003_out_endofpacket;                                                                 // crosser_003:out_endofpacket -> hps_0_h2f_axi_master_agent:read_rp_endofpacket
	wire          crosser_003_out_valid;                                                                       // crosser_003:out_valid -> hps_0_h2f_axi_master_agent:read_rp_valid
	wire          crosser_003_out_startofpacket;                                                               // crosser_003:out_startofpacket -> hps_0_h2f_axi_master_agent:read_rp_startofpacket
	wire  [155:0] crosser_003_out_data;                                                                        // crosser_003:out_data -> hps_0_h2f_axi_master_agent:read_rp_data
	wire    [1:0] crosser_003_out_channel;                                                                     // crosser_003:out_channel -> hps_0_h2f_axi_master_agent:read_rp_channel
	wire          rsp_xbar_demux_src1_endofpacket;                                                             // rsp_xbar_demux:src1_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                   // rsp_xbar_demux:src1_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                           // rsp_xbar_demux:src1_startofpacket -> crosser_003:in_startofpacket
	wire  [155:0] rsp_xbar_demux_src1_data;                                                                    // rsp_xbar_demux:src1_data -> crosser_003:in_data
	wire    [1:0] rsp_xbar_demux_src1_channel;                                                                 // rsp_xbar_demux:src1_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_src1_ready;                                                                   // crosser_003:in_ready -> rsp_xbar_demux:src1_ready

	fpga_sdram_controller_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk               (clk_clk),                                                                  //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                                            //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                                            //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3_emif_0_afi_clk_clk),                                           //          afi_clk.clk
		.afi_half_clk              (),                                                                         //     afi_half_clk.clk
		.afi_reset_n               (mem_if_ddr3_emif_0_afi_reset_reset),                                       //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                                         // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                                                             //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                                                            //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                                                            //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                                          //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                                           //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                                          //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                                            //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                                                         //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                                                         //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                                                          //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                                                       //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                                            //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                                           //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                                         //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                                           //                 .mem_odt
		.avl_ready                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address),            //                 .address
		.avl_rdata_valid           (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata),           //                 .readdata
		.avl_wdata                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata),          //                 .writedata
		.avl_be                    (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable),         //                 .byteenable
		.avl_read_req              (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read),               //                 .read
		.avl_write_req             (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write),              //                 .write
		.avl_size                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount),         //                 .burstcount
		.local_init_done           (),                                                                         //           status.local_init_done
		.local_cal_success         (),                                                                         //                 .local_cal_success
		.local_cal_fail            (),                                                                         //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                                                //              oct.rzqin
		.pll_mem_clk               (),                                                                         //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                                         //                 .pll_write_clk
		.pll_write_clk_pre_phy_clk (),                                                                         //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                                         //                 .pll_addr_cmd_clk
		.pll_locked                (),                                                                         //                 .pll_locked
		.pll_avl_clk               (),                                                                         //                 .pll_avl_clk
		.pll_config_clk            (),                                                                         //                 .pll_config_clk
		.pll_mem_phy_clk           (),                                                                         //                 .pll_mem_phy_clk
		.afi_phy_clk               (),                                                                         //                 .afi_phy_clk
		.pll_avl_phy_clk           ()                                                                          //                 .pll_avl_phy_clk
	);

	fpga_sdram_controller_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps_0 (
		.mem_a       (memory_0_mem_a),               //         memory.mem_a
		.mem_ba      (memory_0_mem_ba),              //               .mem_ba
		.mem_ck      (memory_0_mem_ck),              //               .mem_ck
		.mem_ck_n    (memory_0_mem_ck_n),            //               .mem_ck_n
		.mem_cke     (memory_0_mem_cke),             //               .mem_cke
		.mem_cs_n    (memory_0_mem_cs_n),            //               .mem_cs_n
		.mem_ras_n   (memory_0_mem_ras_n),           //               .mem_ras_n
		.mem_cas_n   (memory_0_mem_cas_n),           //               .mem_cas_n
		.mem_we_n    (memory_0_mem_we_n),            //               .mem_we_n
		.mem_reset_n (memory_0_mem_reset_n),         //               .mem_reset_n
		.mem_dq      (memory_0_mem_dq),              //               .mem_dq
		.mem_dqs     (memory_0_mem_dqs),             //               .mem_dqs
		.mem_dqs_n   (memory_0_mem_dqs_n),           //               .mem_dqs_n
		.mem_odt     (memory_0_mem_odt),             //               .mem_odt
		.mem_dm      (memory_0_mem_dm),              //               .mem_dm
		.oct_rzqin   (memory_0_oct_rzqin),           //               .oct_rzqin
		.h2f_rst_n   (hps_0_h2f_reset_reset),        //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),                      //  h2f_axi_clock.clk
		.h2f_AWID    (hps_0_h2f_axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (hps_0_h2f_axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (hps_0_h2f_axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (hps_0_h2f_axi_master_awsize),  //               .awsize
		.h2f_AWBURST (hps_0_h2f_axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (hps_0_h2f_axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (hps_0_h2f_axi_master_awcache), //               .awcache
		.h2f_AWPROT  (hps_0_h2f_axi_master_awprot),  //               .awprot
		.h2f_AWVALID (hps_0_h2f_axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (hps_0_h2f_axi_master_awready), //               .awready
		.h2f_WID     (hps_0_h2f_axi_master_wid),     //               .wid
		.h2f_WDATA   (hps_0_h2f_axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (hps_0_h2f_axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (hps_0_h2f_axi_master_wlast),   //               .wlast
		.h2f_WVALID  (hps_0_h2f_axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (hps_0_h2f_axi_master_wready),  //               .wready
		.h2f_BID     (hps_0_h2f_axi_master_bid),     //               .bid
		.h2f_BRESP   (hps_0_h2f_axi_master_bresp),   //               .bresp
		.h2f_BVALID  (hps_0_h2f_axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (hps_0_h2f_axi_master_bready),  //               .bready
		.h2f_ARID    (hps_0_h2f_axi_master_arid),    //               .arid
		.h2f_ARADDR  (hps_0_h2f_axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (hps_0_h2f_axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (hps_0_h2f_axi_master_arsize),  //               .arsize
		.h2f_ARBURST (hps_0_h2f_axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (hps_0_h2f_axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (hps_0_h2f_axi_master_arcache), //               .arcache
		.h2f_ARPROT  (hps_0_h2f_axi_master_arprot),  //               .arprot
		.h2f_ARVALID (hps_0_h2f_axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (hps_0_h2f_axi_master_arready), //               .arready
		.h2f_RID     (hps_0_h2f_axi_master_rid),     //               .rid
		.h2f_RDATA   (hps_0_h2f_axi_master_rdata),   //               .rdata
		.h2f_RRESP   (hps_0_h2f_axi_master_rresp),   //               .rresp
		.h2f_RLAST   (hps_0_h2f_axi_master_rlast),   //               .rlast
		.h2f_RVALID  (hps_0_h2f_axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (hps_0_h2f_axi_master_rready)   //               .rready
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (21),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (6),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (30),
		.UAV_BURSTCOUNT_W               (8),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_if_ddr3_emif_0_avl_translator (
		.clk                      (mem_if_ddr3_emif_0_afi_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (12),
		.ADDR_WIDTH                (30),
		.RDATA_WIDTH               (64),
		.WDATA_WIDTH               (64),
		.ADDR_USER_WIDTH           (1),
		.DATA_USER_WIDTH           (1),
		.AXI_BURST_LENGTH_WIDTH    (4),
		.AXI_LOCK_WIDTH            (2),
		.AXI_VERSION               ("AXI3"),
		.WRITE_ISSUING_CAPABILITY  (8),
		.READ_ISSUING_CAPABILITY   (8),
		.PKT_BEGIN_BURST           (131),
		.PKT_CACHE_H               (153),
		.PKT_CACHE_L               (150),
		.PKT_ADDR_SIDEBAND_H       (129),
		.PKT_ADDR_SIDEBAND_L       (129),
		.PKT_PROTECTION_H          (149),
		.PKT_PROTECTION_L          (147),
		.PKT_BURST_SIZE_H          (126),
		.PKT_BURST_SIZE_L          (124),
		.PKT_BURST_TYPE_H          (128),
		.PKT_BURST_TYPE_L          (127),
		.PKT_RESPONSE_STATUS_L     (154),
		.PKT_RESPONSE_STATUS_H     (155),
		.PKT_BURSTWRAP_H           (123),
		.PKT_BURSTWRAP_L           (116),
		.PKT_BYTE_CNT_H            (115),
		.PKT_BYTE_CNT_L            (108),
		.PKT_ADDR_H                (101),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_EXCLUSIVE       (107),
		.PKT_TRANS_LOCK            (106),
		.PKT_TRANS_COMPRESSED_READ (102),
		.PKT_TRANS_POSTED          (103),
		.PKT_TRANS_WRITE           (104),
		.PKT_TRANS_READ            (105),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (133),
		.PKT_SRC_ID_L              (133),
		.PKT_DEST_ID_H             (134),
		.PKT_DEST_ID_L             (134),
		.PKT_THREAD_ID_H           (146),
		.PKT_THREAD_ID_L           (135),
		.PKT_QOS_L                 (132),
		.PKT_QOS_H                 (132),
		.PKT_DATA_SIDEBAND_H       (130),
		.PKT_DATA_SIDEBAND_L       (130),
		.ST_DATA_W                 (156),
		.ST_CHANNEL_W              (2),
		.ID                        (0)
	) hps_0_h2f_axi_master_agent (
		.aclk                   (clk_clk),                                           //              clk.clk
		.aresetn                (~rst_controller_001_reset_out_reset),               //        clk_reset.reset_n
		.write_cp_valid         (hps_0_h2f_axi_master_agent_write_cp_valid),         //         write_cp.valid
		.write_cp_data          (hps_0_h2f_axi_master_agent_write_cp_data),          //                 .data
		.write_cp_startofpacket (hps_0_h2f_axi_master_agent_write_cp_startofpacket), //                 .startofpacket
		.write_cp_endofpacket   (hps_0_h2f_axi_master_agent_write_cp_endofpacket),   //                 .endofpacket
		.write_cp_ready         (hps_0_h2f_axi_master_agent_write_cp_ready),         //                 .ready
		.write_rp_valid         (crosser_002_out_valid),                             //         write_rp.valid
		.write_rp_data          (crosser_002_out_data),                              //                 .data
		.write_rp_channel       (crosser_002_out_channel),                           //                 .channel
		.write_rp_startofpacket (crosser_002_out_startofpacket),                     //                 .startofpacket
		.write_rp_endofpacket   (crosser_002_out_endofpacket),                       //                 .endofpacket
		.write_rp_ready         (crosser_002_out_ready),                             //                 .ready
		.read_cp_valid          (hps_0_h2f_axi_master_agent_read_cp_valid),          //          read_cp.valid
		.read_cp_data           (hps_0_h2f_axi_master_agent_read_cp_data),           //                 .data
		.read_cp_startofpacket  (hps_0_h2f_axi_master_agent_read_cp_startofpacket),  //                 .startofpacket
		.read_cp_endofpacket    (hps_0_h2f_axi_master_agent_read_cp_endofpacket),    //                 .endofpacket
		.read_cp_ready          (hps_0_h2f_axi_master_agent_read_cp_ready),          //                 .ready
		.read_rp_valid          (crosser_003_out_valid),                             //          read_rp.valid
		.read_rp_data           (crosser_003_out_data),                              //                 .data
		.read_rp_channel        (crosser_003_out_channel),                           //                 .channel
		.read_rp_startofpacket  (crosser_003_out_startofpacket),                     //                 .startofpacket
		.read_rp_endofpacket    (crosser_003_out_endofpacket),                       //                 .endofpacket
		.read_rp_ready          (crosser_003_out_ready),                             //                 .ready
		.awid                   (hps_0_h2f_axi_master_awid),                         // altera_axi_slave.awid
		.awaddr                 (hps_0_h2f_axi_master_awaddr),                       //                 .awaddr
		.awlen                  (hps_0_h2f_axi_master_awlen),                        //                 .awlen
		.awsize                 (hps_0_h2f_axi_master_awsize),                       //                 .awsize
		.awburst                (hps_0_h2f_axi_master_awburst),                      //                 .awburst
		.awlock                 (hps_0_h2f_axi_master_awlock),                       //                 .awlock
		.awcache                (hps_0_h2f_axi_master_awcache),                      //                 .awcache
		.awprot                 (hps_0_h2f_axi_master_awprot),                       //                 .awprot
		.awvalid                (hps_0_h2f_axi_master_awvalid),                      //                 .awvalid
		.awready                (hps_0_h2f_axi_master_awready),                      //                 .awready
		.wid                    (hps_0_h2f_axi_master_wid),                          //                 .wid
		.wdata                  (hps_0_h2f_axi_master_wdata),                        //                 .wdata
		.wstrb                  (hps_0_h2f_axi_master_wstrb),                        //                 .wstrb
		.wlast                  (hps_0_h2f_axi_master_wlast),                        //                 .wlast
		.wvalid                 (hps_0_h2f_axi_master_wvalid),                       //                 .wvalid
		.wready                 (hps_0_h2f_axi_master_wready),                       //                 .wready
		.bid                    (hps_0_h2f_axi_master_bid),                          //                 .bid
		.bresp                  (hps_0_h2f_axi_master_bresp),                        //                 .bresp
		.bvalid                 (hps_0_h2f_axi_master_bvalid),                       //                 .bvalid
		.bready                 (hps_0_h2f_axi_master_bready),                       //                 .bready
		.arid                   (hps_0_h2f_axi_master_arid),                         //                 .arid
		.araddr                 (hps_0_h2f_axi_master_araddr),                       //                 .araddr
		.arlen                  (hps_0_h2f_axi_master_arlen),                        //                 .arlen
		.arsize                 (hps_0_h2f_axi_master_arsize),                       //                 .arsize
		.arburst                (hps_0_h2f_axi_master_arburst),                      //                 .arburst
		.arlock                 (hps_0_h2f_axi_master_arlock),                       //                 .arlock
		.arcache                (hps_0_h2f_axi_master_arcache),                      //                 .arcache
		.arprot                 (hps_0_h2f_axi_master_arprot),                       //                 .arprot
		.arvalid                (hps_0_h2f_axi_master_arvalid),                      //                 .arvalid
		.arready                (hps_0_h2f_axi_master_arready),                      //                 .arready
		.rid                    (hps_0_h2f_axi_master_rid),                          //                 .rid
		.rdata                  (hps_0_h2f_axi_master_rdata),                        //                 .rdata
		.rresp                  (hps_0_h2f_axi_master_rresp),                        //                 .rresp
		.rlast                  (hps_0_h2f_axi_master_rlast),                        //                 .rlast
		.rvalid                 (hps_0_h2f_axi_master_rvalid),                       //                 .rvalid
		.rready                 (hps_0_h2f_axi_master_rready),                       //                 .rready
		.awuser                 (1'b0),                                              //      (terminated)
		.aruser                 (1'b0),                                              //      (terminated)
		.awqos                  (4'b0000),                                           //      (terminated)
		.arqos                  (4'b0000),                                           //      (terminated)
		.awregion               (4'b0000),                                           //      (terminated)
		.arregion               (4'b0000),                                           //      (terminated)
		.wuser                  (1'b0),                                              //      (terminated)
		.ruser                  (),                                                  //      (terminated)
		.buser                  ()                                                   //      (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (95),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_SRC_ID_H              (97),
		.PKT_SRC_ID_L              (97),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (98),
		.PKT_BURSTWRAP_H           (87),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (72),
		.PKT_PROTECTION_H          (113),
		.PKT_PROTECTION_L          (111),
		.PKT_RESPONSE_STATUS_H     (119),
		.PKT_RESPONSE_STATUS_L     (118),
		.PKT_BURST_SIZE_H          (90),
		.PKT_BURST_SIZE_L          (88),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (120),
		.AVS_BURSTCOUNT_W          (8),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr3_emif_0_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                 //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                 //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                  //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                           //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                               //                .channel
		.rf_sink_ready           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (121),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr3_emif_0_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2048),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (mem_if_ddr3_emif_0_afi_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	fpga_sdram_controller_addr_router addr_router (
		.sink_ready         (hps_0_h2f_axi_master_agent_write_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_axi_master_agent_write_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_axi_master_agent_write_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_axi_master_agent_write_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_axi_master_agent_write_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                // clk_reset.reset
		.src_ready          (addr_router_src_ready),                             //       src.ready
		.src_valid          (addr_router_src_valid),                             //          .valid
		.src_data           (addr_router_src_data),                              //          .data
		.src_channel        (addr_router_src_channel),                           //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                     //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                        //          .endofpacket
	);

	fpga_sdram_controller_addr_router addr_router_001 (
		.sink_ready         (hps_0_h2f_axi_master_agent_read_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_axi_master_agent_read_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_axi_master_agent_read_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_axi_master_agent_read_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_axi_master_agent_read_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),               // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                        //       src.ready
		.src_valid          (addr_router_001_src_valid),                        //          .valid
		.src_data           (addr_router_001_src_data),                         //          .data
		.src_channel        (addr_router_001_src_channel),                      //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                   //          .endofpacket
	);

	fpga_sdram_controller_id_router id_router (
		.sink_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr3_emif_0_afi_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                               //       src.ready
		.src_valid          (id_router_src_valid),                                                               //          .valid
		.src_data           (id_router_src_data),                                                                //          .data
		.src_channel        (id_router_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                          //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (95),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (72),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (90),
		.PKT_BURST_SIZE_L          (88),
		.PKT_BURST_TYPE_H          (92),
		.PKT_BURST_TYPE_L          (91),
		.PKT_BURSTWRAP_H           (87),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (120),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (79),
		.OUT_BURSTWRAP_H           (87),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter (
		.clk                   (mem_if_ddr3_emif_0_afi_clk_clk),         //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),         // cr0_reset.reset
		.sink0_valid           (width_adapter_cmd_source_valid),         //     sink0.valid
		.sink0_data            (width_adapter_cmd_source_data),          //          .data
		.sink0_channel         (width_adapter_cmd_source_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_cmd_source_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_cmd_source_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_cmd_source_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),            //   source0.valid
		.source0_data          (burst_adapter_source0_data),             //          .data
		.source0_channel       (burst_adapter_source0_channel),          //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket),    //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),      //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)             //          .ready
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (101),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (115),
		.IN_PKT_BYTE_CNT_L             (108),
		.IN_PKT_TRANS_COMPRESSED_READ  (102),
		.IN_PKT_BURSTWRAP_H            (123),
		.IN_PKT_BURSTWRAP_L            (116),
		.IN_PKT_BURST_SIZE_H           (126),
		.IN_PKT_BURST_SIZE_L           (124),
		.IN_PKT_RESPONSE_STATUS_H      (155),
		.IN_PKT_RESPONSE_STATUS_L      (154),
		.IN_PKT_TRANS_EXCLUSIVE        (107),
		.IN_PKT_BURST_TYPE_H           (128),
		.IN_PKT_BURST_TYPE_L           (127),
		.IN_PKT_TRANS_POSTED           (103),
		.IN_ST_DATA_W                  (156),
		.OUT_PKT_ADDR_H                (65),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (72),
		.OUT_PKT_TRANS_COMPRESSED_READ (66),
		.OUT_PKT_TRANS_EXCLUSIVE       (71),
		.OUT_PKT_RESPONSE_STATUS_H     (119),
		.OUT_PKT_RESPONSE_STATUS_L     (118),
		.OUT_PKT_BURST_SIZE_H          (90),
		.OUT_PKT_BURST_SIZE_L          (88),
		.OUT_PKT_BURST_TYPE_H          (92),
		.OUT_PKT_BURST_TYPE_L          (91),
		.OUT_ST_DATA_W                 (120),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (40)
	) width_adapter (
		.clk                   (mem_if_ddr3_emif_0_afi_clk_clk),         //      clock.clk
		.reset                 (rst_controller_reset_out_reset),         //      reset.reset
		.cmd_in_valid          (cmd_xbar_mux_src_valid),                 //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_mux_src_channel),               //           .channel
		.cmd_in_data           (cmd_xbar_mux_src_data),                  //           .data
		.cmd_in_startofpacket  (cmd_xbar_mux_src_startofpacket),         //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_mux_src_endofpacket),           //           .endofpacket
		.cmd_in_ready          (cmd_xbar_mux_src_ready),                 //           .ready
		.cmd_out_ready         (width_adapter_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_src_channel),                  //           .channel
		.rsp_in_data           (id_router_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~mem_if_ddr3_emif_0_afi_reset_reset), // reset_in0.reset
		.clk        (mem_if_ddr3_emif_0_afi_clk_clk),      //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req  (),                                    // (terminated)
		.reset_in1  (1'b0),                                // (terminated)
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	fpga_sdram_controller_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	fpga_sdram_controller_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	fpga_sdram_controller_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (mem_if_ddr3_emif_0_afi_clk_clk), //       clk.clk
		.reset               (rst_controller_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_out_valid),              //          .valid
		.sink0_channel       (crosser_out_channel),            //          .channel
		.sink0_data          (crosser_out_data),               //          .data
		.sink0_startofpacket (crosser_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_001_out_ready),          //     sink1.ready
		.sink1_valid         (crosser_001_out_valid),          //          .valid
		.sink1_channel       (crosser_001_out_channel),        //          .channel
		.sink1_data          (crosser_001_out_data),           //          .data
		.sink1_startofpacket (crosser_001_out_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (crosser_001_out_endofpacket)     //          .endofpacket
	);

	fpga_sdram_controller_rsp_xbar_demux rsp_xbar_demux (
		.clk                (mem_if_ddr3_emif_0_afi_clk_clk),         //       clk.clk
		.reset              (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready         (width_adapter_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),        //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),              //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),              //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),               //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),            //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)         //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (156),
		.BITS_PER_SYMBOL     (156),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (mem_if_ddr3_emif_0_afi_clk_clk),     //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src0_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (156),
		.BITS_PER_SYMBOL     (156),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr3_emif_0_afi_clk_clk),        //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (156),
		.BITS_PER_SYMBOL     (156),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src0_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_002_out_ready),              //           out.ready
		.out_valid         (crosser_002_out_valid),              //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_002_out_channel),            //              .channel
		.out_data          (crosser_002_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (156),
		.BITS_PER_SYMBOL     (156),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src1_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src1_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src1_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src1_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src1_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src1_data),           //              .data
		.out_ready         (crosser_003_out_ready),              //           out.ready
		.out_valid         (crosser_003_out_valid),              //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_003_out_channel),            //              .channel
		.out_data          (crosser_003_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

endmodule
