// fpga_sdram_controller.v

// Generated using ACDS version 13.0sp1 232 at 2015.08.05.16:15:48

`timescale 1 ps / 1 ps
module fpga_sdram_controller (
		input  wire        clk_clk,                            //             clk.clk
		input  wire        reset_reset_n,                      //           reset.reset_n
		output wire [12:0] memory_mem_a,                       //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                      //                .mem_ba
		output wire [0:0]  memory_mem_ck,                      //                .mem_ck
		output wire [0:0]  memory_mem_ck_n,                    //                .mem_ck_n
		output wire [0:0]  memory_mem_cke,                     //                .mem_cke
		output wire [0:0]  memory_mem_cs_n,                    //                .mem_cs_n
		output wire [0:0]  memory_mem_dm,                      //                .mem_dm
		output wire [0:0]  memory_mem_ras_n,                   //                .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                   //                .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                    //                .mem_we_n
		output wire        memory_mem_reset_n,                 //                .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                      //                .mem_dq
		inout  wire [0:0]  memory_mem_dqs,                     //                .mem_dqs
		inout  wire [0:0]  memory_mem_dqs_n,                   //                .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                     //                .mem_odt
		input  wire        oct_rzqin,                          //             oct.rzqin
		output wire        sdram_avl_slave_waitrequest_n,      // sdram_avl_slave.waitrequest_n
		input  wire        sdram_avl_slave_beginbursttransfer, //                .beginbursttransfer
		input  wire [20:0] sdram_avl_slave_address,            //                .address
		output wire        sdram_avl_slave_readdatavalid,      //                .readdatavalid
		output wire [31:0] sdram_avl_slave_readdata,           //                .readdata
		input  wire [31:0] sdram_avl_slave_writedata,          //                .writedata
		input  wire [3:0]  sdram_avl_slave_byteenable,         //                .byteenable
		input  wire        sdram_avl_slave_read,               //                .read
		input  wire        sdram_avl_slave_write,              //                .write
		input  wire [5:0]  sdram_avl_slave_burstcount          //                .burstcount
	);

	fpga_sdram_controller_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk               (clk_clk),                            //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                      //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                      //       soft_reset.reset_n
		.afi_clk                   (),                                   //          afi_clk.clk
		.afi_half_clk              (),                                   //     afi_half_clk.clk
		.afi_reset_n               (),                                   //        afi_reset.reset_n
		.afi_reset_export_n        (),                                   // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                       //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                      //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                      //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                    //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                     //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                    //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                      //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                   //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                   //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                    //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                 //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                      //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                     //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                   //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                     //                 .mem_odt
		.avl_ready                 (sdram_avl_slave_waitrequest_n),      //              avl.waitrequest_n
		.avl_burstbegin            (sdram_avl_slave_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (sdram_avl_slave_address),            //                 .address
		.avl_rdata_valid           (sdram_avl_slave_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (sdram_avl_slave_readdata),           //                 .readdata
		.avl_wdata                 (sdram_avl_slave_writedata),          //                 .writedata
		.avl_be                    (sdram_avl_slave_byteenable),         //                 .byteenable
		.avl_read_req              (sdram_avl_slave_read),               //                 .read
		.avl_write_req             (sdram_avl_slave_write),              //                 .write
		.avl_size                  (sdram_avl_slave_burstcount),         //                 .burstcount
		.local_init_done           (),                                   //           status.local_init_done
		.local_cal_success         (),                                   //                 .local_cal_success
		.local_cal_fail            (),                                   //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                          //              oct.rzqin
		.pll_mem_clk               (),                                   //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                   //                 .pll_write_clk
		.pll_write_clk_pre_phy_clk (),                                   //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                   //                 .pll_addr_cmd_clk
		.pll_locked                (),                                   //                 .pll_locked
		.pll_avl_clk               (),                                   //                 .pll_avl_clk
		.pll_config_clk            (),                                   //                 .pll_config_clk
		.pll_mem_phy_clk           (),                                   //                 .pll_mem_phy_clk
		.afi_phy_clk               (),                                   //                 .afi_phy_clk
		.pll_avl_phy_clk           ()                                    //                 .pll_avl_phy_clk
	);

endmodule
