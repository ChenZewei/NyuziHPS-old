// axi_agent.v

// Generated using ACDS version 13.0sp1 232 at 2015.07.30.10:36:15

`timescale 1 ps / 1 ps
module axi_agent (
		input  wire        clk_clk,            //    clk.clk
		input  wire        reset_reset_n,      //  reset.reset_n
		output wire [12:0] memory_mem_a,       // memory.mem_a
		output wire [2:0]  memory_mem_ba,      //       .mem_ba
		output wire        memory_mem_ck,      //       .mem_ck
		output wire        memory_mem_ck_n,    //       .mem_ck_n
		output wire        memory_mem_cke,     //       .mem_cke
		output wire        memory_mem_cs_n,    //       .mem_cs_n
		output wire        memory_mem_ras_n,   //       .mem_ras_n
		output wire        memory_mem_cas_n,   //       .mem_cas_n
		output wire        memory_mem_we_n,    //       .mem_we_n
		output wire        memory_mem_reset_n, //       .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,      //       .mem_dq
		inout  wire        memory_mem_dqs,     //       .mem_dqs
		inout  wire        memory_mem_dqs_n,   //       .mem_dqs_n
		output wire        memory_mem_odt,     //       .mem_odt
		output wire        memory_mem_dm,      //       .mem_dm
		input  wire        memory_oct_rzqin    //       .oct_rzqin
	);

	wire          hps_0_h2f_axi_master_awvalid;                                            // hps_0:h2f_AWVALID -> id_pad:s0_awvalid
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                             // hps_0:h2f_ARSIZE -> id_pad:s0_arsize
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                             // hps_0:h2f_ARLOCK -> id_pad:s0_arlock
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                            // hps_0:h2f_AWCACHE -> id_pad:s0_awcache
	wire          hps_0_h2f_axi_master_arready;                                            // id_pad:s0_arready -> hps_0:h2f_ARREADY
	wire   [11:0] hps_0_h2f_axi_master_arid;                                               // hps_0:h2f_ARID -> id_pad:s0_arid
	wire          hps_0_h2f_axi_master_rready;                                             // hps_0:h2f_RREADY -> id_pad:s0_rready
	wire          hps_0_h2f_axi_master_bready;                                             // hps_0:h2f_BREADY -> id_pad:s0_bready
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                             // hps_0:h2f_AWSIZE -> id_pad:s0_awsize
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                             // hps_0:h2f_AWPROT -> id_pad:s0_awprot
	wire          hps_0_h2f_axi_master_arvalid;                                            // hps_0:h2f_ARVALID -> id_pad:s0_arvalid
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                             // hps_0:h2f_ARPROT -> id_pad:s0_arprot
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                // id_pad:s0_bid -> hps_0:h2f_BID
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                              // hps_0:h2f_ARLEN -> id_pad:s0_arlen
	wire          hps_0_h2f_axi_master_awready;                                            // id_pad:s0_awready -> hps_0:h2f_AWREADY
	wire   [11:0] hps_0_h2f_axi_master_awid;                                               // hps_0:h2f_AWID -> id_pad:s0_awid
	wire          hps_0_h2f_axi_master_bvalid;                                             // id_pad:s0_bvalid -> hps_0:h2f_BVALID
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                // hps_0:h2f_WID -> id_pad:s0_wid
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                             // hps_0:h2f_AWLOCK -> id_pad:s0_awlock
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                            // hps_0:h2f_AWBURST -> id_pad:s0_awburst
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                              // id_pad:s0_bresp -> hps_0:h2f_BRESP
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                              // hps_0:h2f_WSTRB -> id_pad:s0_wstrb
	wire          hps_0_h2f_axi_master_rvalid;                                             // id_pad:s0_rvalid -> hps_0:h2f_RVALID
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                              // hps_0:h2f_WDATA -> id_pad:s0_wdata
	wire          hps_0_h2f_axi_master_wready;                                             // id_pad:s0_wready -> hps_0:h2f_WREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                            // hps_0:h2f_ARBURST -> id_pad:s0_arburst
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                              // id_pad:s0_rdata -> hps_0:h2f_RDATA
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                             // hps_0:h2f_ARADDR -> id_pad:s0_araddr
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                            // hps_0:h2f_ARCACHE -> id_pad:s0_arcache
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                              // hps_0:h2f_AWLEN -> id_pad:s0_awlen
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                             // hps_0:h2f_AWADDR -> id_pad:s0_awaddr
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                // id_pad:s0_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_wvalid;                                             // hps_0:h2f_WVALID -> id_pad:s0_wvalid
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                              // id_pad:s0_rresp -> hps_0:h2f_RRESP
	wire          hps_0_h2f_axi_master_wlast;                                              // hps_0:h2f_WLAST -> id_pad:s0_wlast
	wire          hps_0_h2f_axi_master_rlast;                                              // id_pad:s0_rlast -> hps_0:h2f_RLAST
	wire          id_pad_m0_awvalid;                                                       // id_pad:m0_awvalid -> id_pad_m0_agent:awvalid
	wire    [2:0] id_pad_m0_arsize;                                                        // id_pad:m0_arsize -> id_pad_m0_agent:arsize
	wire    [1:0] id_pad_m0_arlock;                                                        // id_pad:m0_arlock -> id_pad_m0_agent:arlock
	wire    [3:0] id_pad_m0_awcache;                                                       // id_pad:m0_awcache -> id_pad_m0_agent:awcache
	wire          id_pad_m0_arready;                                                       // id_pad_m0_agent:arready -> id_pad:m0_arready
	wire    [1:0] id_pad_m0_arid;                                                          // id_pad:m0_arid -> id_pad_m0_agent:arid
	wire          id_pad_m0_rready;                                                        // id_pad:m0_rready -> id_pad_m0_agent:rready
	wire          id_pad_m0_bready;                                                        // id_pad:m0_bready -> id_pad_m0_agent:bready
	wire    [2:0] id_pad_m0_awsize;                                                        // id_pad:m0_awsize -> id_pad_m0_agent:awsize
	wire    [2:0] id_pad_m0_awprot;                                                        // id_pad:m0_awprot -> id_pad_m0_agent:awprot
	wire          id_pad_m0_arvalid;                                                       // id_pad:m0_arvalid -> id_pad_m0_agent:arvalid
	wire    [2:0] id_pad_m0_arprot;                                                        // id_pad:m0_arprot -> id_pad_m0_agent:arprot
	wire    [1:0] id_pad_m0_bid;                                                           // id_pad_m0_agent:bid -> id_pad:m0_bid
	wire    [3:0] id_pad_m0_arlen;                                                         // id_pad:m0_arlen -> id_pad_m0_agent:arlen
	wire          id_pad_m0_awready;                                                       // id_pad_m0_agent:awready -> id_pad:m0_awready
	wire    [1:0] id_pad_m0_awid;                                                          // id_pad:m0_awid -> id_pad_m0_agent:awid
	wire          id_pad_m0_bvalid;                                                        // id_pad_m0_agent:bvalid -> id_pad:m0_bvalid
	wire    [1:0] id_pad_m0_wid;                                                           // id_pad:m0_wid -> id_pad_m0_agent:wid
	wire    [1:0] id_pad_m0_awlock;                                                        // id_pad:m0_awlock -> id_pad_m0_agent:awlock
	wire    [1:0] id_pad_m0_awburst;                                                       // id_pad:m0_awburst -> id_pad_m0_agent:awburst
	wire    [1:0] id_pad_m0_bresp;                                                         // id_pad_m0_agent:bresp -> id_pad:m0_bresp
	wire    [4:0] id_pad_m0_aruser;                                                        // id_pad:m0_aruser -> id_pad_m0_agent:aruser
	wire    [4:0] id_pad_m0_awuser;                                                        // id_pad:m0_awuser -> id_pad_m0_agent:awuser
	wire    [7:0] id_pad_m0_wstrb;                                                         // id_pad:m0_wstrb -> id_pad_m0_agent:wstrb
	wire          id_pad_m0_rvalid;                                                        // id_pad_m0_agent:rvalid -> id_pad:m0_rvalid
	wire    [1:0] id_pad_m0_arburst;                                                       // id_pad:m0_arburst -> id_pad_m0_agent:arburst
	wire   [63:0] id_pad_m0_wdata;                                                         // id_pad:m0_wdata -> id_pad_m0_agent:wdata
	wire          id_pad_m0_wready;                                                        // id_pad_m0_agent:wready -> id_pad:m0_wready
	wire   [63:0] id_pad_m0_rdata;                                                         // id_pad_m0_agent:rdata -> id_pad:m0_rdata
	wire   [29:0] id_pad_m0_araddr;                                                        // id_pad:m0_araddr -> id_pad_m0_agent:araddr
	wire    [3:0] id_pad_m0_arcache;                                                       // id_pad:m0_arcache -> id_pad_m0_agent:arcache
	wire    [3:0] id_pad_m0_awlen;                                                         // id_pad:m0_awlen -> id_pad_m0_agent:awlen
	wire   [29:0] id_pad_m0_awaddr;                                                        // id_pad:m0_awaddr -> id_pad_m0_agent:awaddr
	wire    [1:0] id_pad_m0_rid;                                                           // id_pad_m0_agent:rid -> id_pad:m0_rid
	wire          id_pad_m0_wvalid;                                                        // id_pad:m0_wvalid -> id_pad_m0_agent:wvalid
	wire    [1:0] id_pad_m0_rresp;                                                         // id_pad_m0_agent:rresp -> id_pad:m0_rresp
	wire          id_pad_m0_wlast;                                                         // id_pad:m0_wlast -> id_pad_m0_agent:wlast
	wire          id_pad_m0_rlast;                                                         // id_pad_m0_agent:rlast -> id_pad:m0_rlast
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awvalid; // merlin_axi_master_ni_0_altera_axi_slave_agent:awvalid -> merlin_axi_master_ni_0:awvalid
	wire    [2:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arsize;  // merlin_axi_master_ni_0_altera_axi_slave_agent:arsize -> merlin_axi_master_ni_0:arsize
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlock;  // merlin_axi_master_ni_0_altera_axi_slave_agent:arlock -> merlin_axi_master_ni_0:arlock
	wire    [3:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awcache; // merlin_axi_master_ni_0_altera_axi_slave_agent:awcache -> merlin_axi_master_ni_0:awcache
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arready; // merlin_axi_master_ni_0:arready -> merlin_axi_master_ni_0_altera_axi_slave_agent:arready
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arid;    // merlin_axi_master_ni_0_altera_axi_slave_agent:arid -> merlin_axi_master_ni_0:arid
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rready;  // merlin_axi_master_ni_0_altera_axi_slave_agent:rready -> merlin_axi_master_ni_0:rready
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bready;  // merlin_axi_master_ni_0_altera_axi_slave_agent:bready -> merlin_axi_master_ni_0:bready
	wire    [2:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awsize;  // merlin_axi_master_ni_0_altera_axi_slave_agent:awsize -> merlin_axi_master_ni_0:awsize
	wire    [2:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awprot;  // merlin_axi_master_ni_0_altera_axi_slave_agent:awprot -> merlin_axi_master_ni_0:awprot
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arvalid; // merlin_axi_master_ni_0_altera_axi_slave_agent:arvalid -> merlin_axi_master_ni_0:arvalid
	wire    [2:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arprot;  // merlin_axi_master_ni_0_altera_axi_slave_agent:arprot -> merlin_axi_master_ni_0:arprot
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bid;     // merlin_axi_master_ni_0:bid -> merlin_axi_master_ni_0_altera_axi_slave_agent:bid
	wire    [3:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlen;   // merlin_axi_master_ni_0_altera_axi_slave_agent:arlen -> merlin_axi_master_ni_0:arlen
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awready; // merlin_axi_master_ni_0:awready -> merlin_axi_master_ni_0_altera_axi_slave_agent:awready
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awid;    // merlin_axi_master_ni_0_altera_axi_slave_agent:awid -> merlin_axi_master_ni_0:awid
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bvalid;  // merlin_axi_master_ni_0:bvalid -> merlin_axi_master_ni_0_altera_axi_slave_agent:bvalid
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wid;     // merlin_axi_master_ni_0_altera_axi_slave_agent:wid -> merlin_axi_master_ni_0:wid
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlock;  // merlin_axi_master_ni_0_altera_axi_slave_agent:awlock -> merlin_axi_master_ni_0:awlock
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awburst; // merlin_axi_master_ni_0_altera_axi_slave_agent:awburst -> merlin_axi_master_ni_0:awburst
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bresp;   // merlin_axi_master_ni_0:bresp -> merlin_axi_master_ni_0_altera_axi_slave_agent:bresp
	wire    [4:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_aruser;  // merlin_axi_master_ni_0_altera_axi_slave_agent:aruser -> merlin_axi_master_ni_0:aruser
	wire    [4:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awuser;  // merlin_axi_master_ni_0_altera_axi_slave_agent:awuser -> merlin_axi_master_ni_0:awuser
	wire    [3:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wstrb;   // merlin_axi_master_ni_0_altera_axi_slave_agent:wstrb -> merlin_axi_master_ni_0:wstrb
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rvalid;  // merlin_axi_master_ni_0:rvalid -> merlin_axi_master_ni_0_altera_axi_slave_agent:rvalid
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arburst; // merlin_axi_master_ni_0_altera_axi_slave_agent:arburst -> merlin_axi_master_ni_0:arburst
	wire   [31:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wdata;   // merlin_axi_master_ni_0_altera_axi_slave_agent:wdata -> merlin_axi_master_ni_0:wdata
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wready;  // merlin_axi_master_ni_0:wready -> merlin_axi_master_ni_0_altera_axi_slave_agent:wready
	wire   [31:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rdata;   // merlin_axi_master_ni_0:rdata -> merlin_axi_master_ni_0_altera_axi_slave_agent:rdata
	wire   [29:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_araddr;  // merlin_axi_master_ni_0_altera_axi_slave_agent:araddr -> merlin_axi_master_ni_0:araddr
	wire    [3:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arcache; // merlin_axi_master_ni_0_altera_axi_slave_agent:arcache -> merlin_axi_master_ni_0:arcache
	wire    [3:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlen;   // merlin_axi_master_ni_0_altera_axi_slave_agent:awlen -> merlin_axi_master_ni_0:awlen
	wire   [29:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awaddr;  // merlin_axi_master_ni_0_altera_axi_slave_agent:awaddr -> merlin_axi_master_ni_0:awaddr
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rid;     // merlin_axi_master_ni_0:rid -> merlin_axi_master_ni_0_altera_axi_slave_agent:rid
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wvalid;  // merlin_axi_master_ni_0_altera_axi_slave_agent:wvalid -> merlin_axi_master_ni_0:wvalid
	wire    [1:0] merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rresp;   // merlin_axi_master_ni_0:rresp -> merlin_axi_master_ni_0_altera_axi_slave_agent:rresp
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wlast;   // merlin_axi_master_ni_0_altera_axi_slave_agent:wlast -> merlin_axi_master_ni_0:wlast
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rlast;   // merlin_axi_master_ni_0:rlast -> merlin_axi_master_ni_0_altera_axi_slave_agent:rlast
	wire          id_pad_m0_agent_write_cp_endofpacket;                                    // id_pad_m0_agent:write_cp_endofpacket -> addr_router:sink_endofpacket
	wire          id_pad_m0_agent_write_cp_valid;                                          // id_pad_m0_agent:write_cp_valid -> addr_router:sink_valid
	wire          id_pad_m0_agent_write_cp_startofpacket;                                  // id_pad_m0_agent:write_cp_startofpacket -> addr_router:sink_startofpacket
	wire  [149:0] id_pad_m0_agent_write_cp_data;                                           // id_pad_m0_agent:write_cp_data -> addr_router:sink_data
	wire          id_pad_m0_agent_write_cp_ready;                                          // addr_router:sink_ready -> id_pad_m0_agent:write_cp_ready
	wire          id_pad_m0_agent_read_cp_endofpacket;                                     // id_pad_m0_agent:read_cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          id_pad_m0_agent_read_cp_valid;                                           // id_pad_m0_agent:read_cp_valid -> addr_router_001:sink_valid
	wire          id_pad_m0_agent_read_cp_startofpacket;                                   // id_pad_m0_agent:read_cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [149:0] id_pad_m0_agent_read_cp_data;                                            // id_pad_m0_agent:read_cp_data -> addr_router_001:sink_data
	wire          id_pad_m0_agent_read_cp_ready;                                           // addr_router_001:sink_ready -> id_pad_m0_agent:read_cp_ready
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_endofpacket;      // merlin_axi_master_ni_0_altera_axi_slave_agent:write_rp_endofpacket -> id_router:sink_endofpacket
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_valid;            // merlin_axi_master_ni_0_altera_axi_slave_agent:write_rp_valid -> id_router:sink_valid
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_startofpacket;    // merlin_axi_master_ni_0_altera_axi_slave_agent:write_rp_startofpacket -> id_router:sink_startofpacket
	wire  [113:0] merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_data;             // merlin_axi_master_ni_0_altera_axi_slave_agent:write_rp_data -> id_router:sink_data
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_ready;            // id_router:sink_ready -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_rp_ready
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_endofpacket;       // merlin_axi_master_ni_0_altera_axi_slave_agent:read_rp_endofpacket -> id_router_001:sink_endofpacket
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_valid;             // merlin_axi_master_ni_0_altera_axi_slave_agent:read_rp_valid -> id_router_001:sink_valid
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_startofpacket;     // merlin_axi_master_ni_0_altera_axi_slave_agent:read_rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [113:0] merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_data;              // merlin_axi_master_ni_0_altera_axi_slave_agent:read_rp_data -> id_router_001:sink_data
	wire          merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_ready;             // id_router_001:sink_ready -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_rp_ready
	wire          burst_adapter_source0_endofpacket;                                       // burst_adapter:source0_endofpacket -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_endofpacket
	wire          burst_adapter_source0_valid;                                             // burst_adapter:source0_valid -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_valid
	wire          burst_adapter_source0_startofpacket;                                     // burst_adapter:source0_startofpacket -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_startofpacket
	wire  [113:0] burst_adapter_source0_data;                                              // burst_adapter:source0_data -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_data
	wire          burst_adapter_source0_ready;                                             // merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                           // burst_adapter:source0_channel -> merlin_axi_master_ni_0_altera_axi_slave_agent:write_cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                   // burst_adapter_001:source0_endofpacket -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                         // burst_adapter_001:source0_valid -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                 // burst_adapter_001:source0_startofpacket -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_startofpacket
	wire  [113:0] burst_adapter_001_source0_data;                                          // burst_adapter_001:source0_data -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_data
	wire          burst_adapter_001_source0_ready;                                         // merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_ready -> burst_adapter_001:source0_ready
	wire    [1:0] burst_adapter_001_source0_channel;                                       // burst_adapter_001:source0_channel -> merlin_axi_master_ni_0_altera_axi_slave_agent:read_cp_channel
	wire          width_adapter_cmd_source_endofpacket;                                    // width_adapter:cmd_out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_cmd_source_valid;                                          // width_adapter:cmd_out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_cmd_source_startofpacket;                                  // width_adapter:cmd_out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [113:0] width_adapter_cmd_source_data;                                           // width_adapter:cmd_out_data -> burst_adapter:sink0_data
	wire    [1:0] width_adapter_cmd_source_channel;                                        // width_adapter:cmd_out_channel -> burst_adapter:sink0_channel
	wire          width_adapter_cmd_source_ready;                                          // burst_adapter:sink0_ready -> width_adapter:cmd_out_ready
	wire          id_router_src_endofpacket;                                               // id_router:src_endofpacket -> width_adapter:rsp_in_endofpacket
	wire          id_router_src_valid;                                                     // id_router:src_valid -> width_adapter:rsp_in_valid
	wire          id_router_src_startofpacket;                                             // id_router:src_startofpacket -> width_adapter:rsp_in_startofpacket
	wire  [113:0] id_router_src_data;                                                      // id_router:src_data -> width_adapter:rsp_in_data
	wire    [1:0] id_router_src_channel;                                                   // id_router:src_channel -> width_adapter:rsp_in_channel
	wire          id_router_src_ready;                                                     // width_adapter:rsp_in_ready -> id_router:src_ready
	wire          width_adapter_001_cmd_source_endofpacket;                                // width_adapter_001:cmd_out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_001_cmd_source_valid;                                      // width_adapter_001:cmd_out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_001_cmd_source_startofpacket;                              // width_adapter_001:cmd_out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [113:0] width_adapter_001_cmd_source_data;                                       // width_adapter_001:cmd_out_data -> burst_adapter_001:sink0_data
	wire    [1:0] width_adapter_001_cmd_source_channel;                                    // width_adapter_001:cmd_out_channel -> burst_adapter_001:sink0_channel
	wire          width_adapter_001_cmd_source_ready;                                      // burst_adapter_001:sink0_ready -> width_adapter_001:cmd_out_ready
	wire          id_router_001_src_endofpacket;                                           // id_router_001:src_endofpacket -> width_adapter_001:rsp_in_endofpacket
	wire          id_router_001_src_valid;                                                 // id_router_001:src_valid -> width_adapter_001:rsp_in_valid
	wire          id_router_001_src_startofpacket;                                         // id_router_001:src_startofpacket -> width_adapter_001:rsp_in_startofpacket
	wire  [113:0] id_router_001_src_data;                                                  // id_router_001:src_data -> width_adapter_001:rsp_in_data
	wire    [1:0] id_router_001_src_channel;                                               // id_router_001:src_channel -> width_adapter_001:rsp_in_channel
	wire          id_router_001_src_ready;                                                 // width_adapter_001:rsp_in_ready -> id_router_001:src_ready
	wire          rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, id_pad:aresetn, id_pad_m0_agent:aresetn, id_router:reset, id_router_001:reset, merlin_axi_master_ni_0:aresetn, merlin_axi_master_ni_0_altera_axi_slave_agent:aresetn, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, width_adapter:reset, width_adapter_001:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                         // cmd_xbar_demux:src0_endofpacket -> width_adapter:cmd_in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                               // cmd_xbar_demux:src0_valid -> width_adapter:cmd_in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                       // cmd_xbar_demux:src0_startofpacket -> width_adapter:cmd_in_startofpacket
	wire  [149:0] cmd_xbar_demux_src0_data;                                                // cmd_xbar_demux:src0_data -> width_adapter:cmd_in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                             // cmd_xbar_demux:src0_channel -> width_adapter:cmd_in_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                     // cmd_xbar_demux_001:src0_endofpacket -> width_adapter_001:cmd_in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                           // cmd_xbar_demux_001:src0_valid -> width_adapter_001:cmd_in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                   // cmd_xbar_demux_001:src0_startofpacket -> width_adapter_001:cmd_in_startofpacket
	wire  [149:0] cmd_xbar_demux_001_src0_data;                                            // cmd_xbar_demux_001:src0_data -> width_adapter_001:cmd_in_data
	wire    [1:0] cmd_xbar_demux_001_src0_channel;                                         // cmd_xbar_demux_001:src0_channel -> width_adapter_001:cmd_in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                         // rsp_xbar_demux:src0_endofpacket -> id_pad_m0_agent:write_rp_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                               // rsp_xbar_demux:src0_valid -> id_pad_m0_agent:write_rp_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                       // rsp_xbar_demux:src0_startofpacket -> id_pad_m0_agent:write_rp_startofpacket
	wire  [149:0] rsp_xbar_demux_src0_data;                                                // rsp_xbar_demux:src0_data -> id_pad_m0_agent:write_rp_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                             // rsp_xbar_demux:src0_channel -> id_pad_m0_agent:write_rp_channel
	wire          rsp_xbar_demux_001_src0_endofpacket;                                     // rsp_xbar_demux_001:src0_endofpacket -> id_pad_m0_agent:read_rp_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                           // rsp_xbar_demux_001:src0_valid -> id_pad_m0_agent:read_rp_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                   // rsp_xbar_demux_001:src0_startofpacket -> id_pad_m0_agent:read_rp_startofpacket
	wire  [149:0] rsp_xbar_demux_001_src0_data;                                            // rsp_xbar_demux_001:src0_data -> id_pad_m0_agent:read_rp_data
	wire    [1:0] rsp_xbar_demux_001_src0_channel;                                         // rsp_xbar_demux_001:src0_channel -> id_pad_m0_agent:read_rp_channel
	wire          addr_router_src_endofpacket;                                             // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                   // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                           // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [149:0] addr_router_src_data;                                                    // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] addr_router_src_channel;                                                 // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                   // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_demux_src0_ready;                                               // id_pad_m0_agent:write_rp_ready -> rsp_xbar_demux:src0_ready
	wire          addr_router_001_src_endofpacket;                                         // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                               // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                       // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [149:0] addr_router_001_src_data;                                                // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [1:0] addr_router_001_src_channel;                                             // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                               // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_demux_001_src0_ready;                                           // id_pad_m0_agent:read_rp_ready -> rsp_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_src0_ready;                                               // width_adapter:cmd_in_ready -> cmd_xbar_demux:src0_ready
	wire          width_adapter_rsp_source_endofpacket;                                    // width_adapter:rsp_out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_rsp_source_valid;                                          // width_adapter:rsp_out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_rsp_source_startofpacket;                                  // width_adapter:rsp_out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [149:0] width_adapter_rsp_source_data;                                           // width_adapter:rsp_out_data -> rsp_xbar_demux:sink_data
	wire    [1:0] width_adapter_rsp_source_channel;                                        // width_adapter:rsp_out_channel -> rsp_xbar_demux:sink_channel
	wire          width_adapter_rsp_source_ready;                                          // rsp_xbar_demux:sink_ready -> width_adapter:rsp_out_ready
	wire          cmd_xbar_demux_001_src0_ready;                                           // width_adapter_001:cmd_in_ready -> cmd_xbar_demux_001:src0_ready
	wire          width_adapter_001_rsp_source_endofpacket;                                // width_adapter_001:rsp_out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_rsp_source_valid;                                      // width_adapter_001:rsp_out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_rsp_source_startofpacket;                              // width_adapter_001:rsp_out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [149:0] width_adapter_001_rsp_source_data;                                       // width_adapter_001:rsp_out_data -> rsp_xbar_demux_001:sink_data
	wire    [1:0] width_adapter_001_rsp_source_channel;                                    // width_adapter_001:rsp_out_channel -> rsp_xbar_demux_001:sink_channel
	wire          width_adapter_001_rsp_source_ready;                                      // rsp_xbar_demux_001:sink_ready -> width_adapter_001:rsp_out_ready

	axi_agent_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.mem_a          (memory_mem_a),                 //            memory.mem_a
		.mem_ba         (memory_mem_ba),                //                  .mem_ba
		.mem_ck         (memory_mem_ck),                //                  .mem_ck
		.mem_ck_n       (memory_mem_ck_n),              //                  .mem_ck_n
		.mem_cke        (memory_mem_cke),               //                  .mem_cke
		.mem_cs_n       (memory_mem_cs_n),              //                  .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),             //                  .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),             //                  .mem_cas_n
		.mem_we_n       (memory_mem_we_n),              //                  .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),           //                  .mem_reset_n
		.mem_dq         (memory_mem_dq),                //                  .mem_dq
		.mem_dqs        (memory_mem_dqs),               //                  .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),             //                  .mem_dqs_n
		.mem_odt        (memory_mem_odt),               //                  .mem_odt
		.mem_dm         (memory_mem_dm),                //                  .mem_dm
		.oct_rzqin      (memory_oct_rzqin),             //                  .oct_rzqin
		.h2f_rst_n      (),                             //         h2f_reset.reset_n
		.h2f_axi_clk    (clk_clk),                      //     h2f_axi_clock.clk
		.h2f_AWID       (hps_0_h2f_axi_master_awid),    //    h2f_axi_master.awid
		.h2f_AWADDR     (hps_0_h2f_axi_master_awaddr),  //                  .awaddr
		.h2f_AWLEN      (hps_0_h2f_axi_master_awlen),   //                  .awlen
		.h2f_AWSIZE     (hps_0_h2f_axi_master_awsize),  //                  .awsize
		.h2f_AWBURST    (hps_0_h2f_axi_master_awburst), //                  .awburst
		.h2f_AWLOCK     (hps_0_h2f_axi_master_awlock),  //                  .awlock
		.h2f_AWCACHE    (hps_0_h2f_axi_master_awcache), //                  .awcache
		.h2f_AWPROT     (hps_0_h2f_axi_master_awprot),  //                  .awprot
		.h2f_AWVALID    (hps_0_h2f_axi_master_awvalid), //                  .awvalid
		.h2f_AWREADY    (hps_0_h2f_axi_master_awready), //                  .awready
		.h2f_WID        (hps_0_h2f_axi_master_wid),     //                  .wid
		.h2f_WDATA      (hps_0_h2f_axi_master_wdata),   //                  .wdata
		.h2f_WSTRB      (hps_0_h2f_axi_master_wstrb),   //                  .wstrb
		.h2f_WLAST      (hps_0_h2f_axi_master_wlast),   //                  .wlast
		.h2f_WVALID     (hps_0_h2f_axi_master_wvalid),  //                  .wvalid
		.h2f_WREADY     (hps_0_h2f_axi_master_wready),  //                  .wready
		.h2f_BID        (hps_0_h2f_axi_master_bid),     //                  .bid
		.h2f_BRESP      (hps_0_h2f_axi_master_bresp),   //                  .bresp
		.h2f_BVALID     (hps_0_h2f_axi_master_bvalid),  //                  .bvalid
		.h2f_BREADY     (hps_0_h2f_axi_master_bready),  //                  .bready
		.h2f_ARID       (hps_0_h2f_axi_master_arid),    //                  .arid
		.h2f_ARADDR     (hps_0_h2f_axi_master_araddr),  //                  .araddr
		.h2f_ARLEN      (hps_0_h2f_axi_master_arlen),   //                  .arlen
		.h2f_ARSIZE     (hps_0_h2f_axi_master_arsize),  //                  .arsize
		.h2f_ARBURST    (hps_0_h2f_axi_master_arburst), //                  .arburst
		.h2f_ARLOCK     (hps_0_h2f_axi_master_arlock),  //                  .arlock
		.h2f_ARCACHE    (hps_0_h2f_axi_master_arcache), //                  .arcache
		.h2f_ARPROT     (hps_0_h2f_axi_master_arprot),  //                  .arprot
		.h2f_ARVALID    (hps_0_h2f_axi_master_arvalid), //                  .arvalid
		.h2f_ARREADY    (hps_0_h2f_axi_master_arready), //                  .arready
		.h2f_RID        (hps_0_h2f_axi_master_rid),     //                  .rid
		.h2f_RDATA      (hps_0_h2f_axi_master_rdata),   //                  .rdata
		.h2f_RRESP      (hps_0_h2f_axi_master_rresp),   //                  .rresp
		.h2f_RLAST      (hps_0_h2f_axi_master_rlast),   //                  .rlast
		.h2f_RVALID     (hps_0_h2f_axi_master_rvalid),  //                  .rvalid
		.h2f_RREADY     (hps_0_h2f_axi_master_rready),  //                  .rready
		.f2h_axi_clk    (clk_clk),                      //     f2h_axi_clock.clk
		.f2h_AWID       (),                             //     f2h_axi_slave.awid
		.f2h_AWADDR     (),                             //                  .awaddr
		.f2h_AWLEN      (),                             //                  .awlen
		.f2h_AWSIZE     (),                             //                  .awsize
		.f2h_AWBURST    (),                             //                  .awburst
		.f2h_AWLOCK     (),                             //                  .awlock
		.f2h_AWCACHE    (),                             //                  .awcache
		.f2h_AWPROT     (),                             //                  .awprot
		.f2h_AWVALID    (),                             //                  .awvalid
		.f2h_AWREADY    (),                             //                  .awready
		.f2h_AWUSER     (),                             //                  .awuser
		.f2h_WID        (),                             //                  .wid
		.f2h_WDATA      (),                             //                  .wdata
		.f2h_WSTRB      (),                             //                  .wstrb
		.f2h_WLAST      (),                             //                  .wlast
		.f2h_WVALID     (),                             //                  .wvalid
		.f2h_WREADY     (),                             //                  .wready
		.f2h_BID        (),                             //                  .bid
		.f2h_BRESP      (),                             //                  .bresp
		.f2h_BVALID     (),                             //                  .bvalid
		.f2h_BREADY     (),                             //                  .bready
		.f2h_ARID       (),                             //                  .arid
		.f2h_ARADDR     (),                             //                  .araddr
		.f2h_ARLEN      (),                             //                  .arlen
		.f2h_ARSIZE     (),                             //                  .arsize
		.f2h_ARBURST    (),                             //                  .arburst
		.f2h_ARLOCK     (),                             //                  .arlock
		.f2h_ARCACHE    (),                             //                  .arcache
		.f2h_ARPROT     (),                             //                  .arprot
		.f2h_ARVALID    (),                             //                  .arvalid
		.f2h_ARREADY    (),                             //                  .arready
		.f2h_ARUSER     (),                             //                  .aruser
		.f2h_RID        (),                             //                  .rid
		.f2h_RDATA      (),                             //                  .rdata
		.f2h_RRESP      (),                             //                  .rresp
		.f2h_RLAST      (),                             //                  .rlast
		.f2h_RVALID     (),                             //                  .rvalid
		.f2h_RREADY     (),                             //                  .rready
		.h2f_lw_axi_clk (clk_clk),                      //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (),                             // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (),                             //                  .awaddr
		.h2f_lw_AWLEN   (),                             //                  .awlen
		.h2f_lw_AWSIZE  (),                             //                  .awsize
		.h2f_lw_AWBURST (),                             //                  .awburst
		.h2f_lw_AWLOCK  (),                             //                  .awlock
		.h2f_lw_AWCACHE (),                             //                  .awcache
		.h2f_lw_AWPROT  (),                             //                  .awprot
		.h2f_lw_AWVALID (),                             //                  .awvalid
		.h2f_lw_AWREADY (),                             //                  .awready
		.h2f_lw_WID     (),                             //                  .wid
		.h2f_lw_WDATA   (),                             //                  .wdata
		.h2f_lw_WSTRB   (),                             //                  .wstrb
		.h2f_lw_WLAST   (),                             //                  .wlast
		.h2f_lw_WVALID  (),                             //                  .wvalid
		.h2f_lw_WREADY  (),                             //                  .wready
		.h2f_lw_BID     (),                             //                  .bid
		.h2f_lw_BRESP   (),                             //                  .bresp
		.h2f_lw_BVALID  (),                             //                  .bvalid
		.h2f_lw_BREADY  (),                             //                  .bready
		.h2f_lw_ARID    (),                             //                  .arid
		.h2f_lw_ARADDR  (),                             //                  .araddr
		.h2f_lw_ARLEN   (),                             //                  .arlen
		.h2f_lw_ARSIZE  (),                             //                  .arsize
		.h2f_lw_ARBURST (),                             //                  .arburst
		.h2f_lw_ARLOCK  (),                             //                  .arlock
		.h2f_lw_ARCACHE (),                             //                  .arcache
		.h2f_lw_ARPROT  (),                             //                  .arprot
		.h2f_lw_ARVALID (),                             //                  .arvalid
		.h2f_lw_ARREADY (),                             //                  .arready
		.h2f_lw_RID     (),                             //                  .rid
		.h2f_lw_RDATA   (),                             //                  .rdata
		.h2f_lw_RRESP   (),                             //                  .rresp
		.h2f_lw_RLAST   (),                             //                  .rlast
		.h2f_lw_RVALID  (),                             //                  .rvalid
		.h2f_lw_RREADY  ()                              //                  .rready
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (2),
		.ADDR_WIDTH                (30),
		.RDATA_WIDTH               (32),
		.WDATA_WIDTH               (32),
		.ADDR_USER_WIDTH           (5),
		.DATA_USER_WIDTH           (8),
		.AXI_BURST_LENGTH_WIDTH    (4),
		.AXI_LOCK_WIDTH            (2),
		.AXI_VERSION               ("AXI3"),
		.WRITE_ISSUING_CAPABILITY  (16),
		.READ_ISSUING_CAPABILITY   (16),
		.PKT_BEGIN_BURST           (104),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_ADDR_SIDEBAND_H       (99),
		.PKT_ADDR_SIDEBAND_L       (92),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (73),
		.PKT_ADDR_L                (42),
		.PKT_TRANS_EXCLUSIVE       (81),
		.PKT_TRANS_LOCK            (105),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (40),
		.PKT_TRANS_WRITE           (39),
		.PKT_TRANS_READ            (38),
		.PKT_DATA_H                (37),
		.PKT_DATA_L                (6),
		.PKT_BYTEEN_H              (5),
		.PKT_BYTEEN_L              (2),
		.PKT_SRC_ID_H              (1),
		.PKT_SRC_ID_L              (1),
		.PKT_DEST_ID_H             (0),
		.PKT_DEST_ID_L             (0),
		.PKT_THREAD_ID_H           (109),
		.PKT_THREAD_ID_L           (108),
		.PKT_QOS_L                 (110),
		.PKT_QOS_H                 (113),
		.PKT_DATA_SIDEBAND_H       (121),
		.PKT_DATA_SIDEBAND_L       (114),
		.ST_DATA_W                 (122),
		.ST_CHANNEL_W              (1),
		.ID                        (1)
	) merlin_axi_master_ni_0 (
		.aclk                   (clk_clk),                                                                 //              clk.clk
		.aresetn                (~rst_controller_reset_out_reset),                                         //        clk_reset.reset_n
		.write_cp_valid         (),                                                                        //         write_cp.valid
		.write_cp_data          (),                                                                        //                 .data
		.write_cp_startofpacket (),                                                                        //                 .startofpacket
		.write_cp_endofpacket   (),                                                                        //                 .endofpacket
		.write_cp_ready         (),                                                                        //                 .ready
		.write_rp_valid         (),                                                                        //         write_rp.valid
		.write_rp_data          (),                                                                        //                 .data
		.write_rp_channel       (),                                                                        //                 .channel
		.write_rp_startofpacket (),                                                                        //                 .startofpacket
		.write_rp_endofpacket   (),                                                                        //                 .endofpacket
		.write_rp_ready         (),                                                                        //                 .ready
		.read_cp_valid          (),                                                                        //          read_cp.valid
		.read_cp_data           (),                                                                        //                 .data
		.read_cp_startofpacket  (),                                                                        //                 .startofpacket
		.read_cp_endofpacket    (),                                                                        //                 .endofpacket
		.read_cp_ready          (),                                                                        //                 .ready
		.read_rp_valid          (),                                                                        //          read_rp.valid
		.read_rp_data           (),                                                                        //                 .data
		.read_rp_channel        (),                                                                        //                 .channel
		.read_rp_startofpacket  (),                                                                        //                 .startofpacket
		.read_rp_endofpacket    (),                                                                        //                 .endofpacket
		.read_rp_ready          (),                                                                        //                 .ready
		.awid                   (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awid),    // altera_axi_slave.awid
		.awaddr                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awaddr),  //                 .awaddr
		.awlen                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlen),   //                 .awlen
		.awsize                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awsize),  //                 .awsize
		.awburst                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awburst), //                 .awburst
		.awlock                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlock),  //                 .awlock
		.awcache                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awcache), //                 .awcache
		.awprot                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awprot),  //                 .awprot
		.awuser                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awuser),  //                 .awuser
		.awvalid                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awvalid), //                 .awvalid
		.awready                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awready), //                 .awready
		.wid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wid),     //                 .wid
		.wdata                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wdata),   //                 .wdata
		.wstrb                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wstrb),   //                 .wstrb
		.wlast                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wlast),   //                 .wlast
		.wvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wvalid),  //                 .wvalid
		.wready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wready),  //                 .wready
		.bid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bid),     //                 .bid
		.bresp                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bresp),   //                 .bresp
		.bvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bvalid),  //                 .bvalid
		.bready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bready),  //                 .bready
		.arid                   (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arid),    //                 .arid
		.araddr                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_araddr),  //                 .araddr
		.arlen                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlen),   //                 .arlen
		.arsize                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arsize),  //                 .arsize
		.arburst                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arburst), //                 .arburst
		.arlock                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlock),  //                 .arlock
		.arcache                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arcache), //                 .arcache
		.arprot                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arprot),  //                 .arprot
		.aruser                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_aruser),  //                 .aruser
		.arvalid                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arvalid), //                 .arvalid
		.arready                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arready), //                 .arready
		.rid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rid),     //                 .rid
		.rdata                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rdata),   //                 .rdata
		.rresp                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rresp),   //                 .rresp
		.rlast                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rlast),   //                 .rlast
		.rvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rvalid),  //                 .rvalid
		.rready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rready),  //                 .rready
		.awqos                  (4'b0000),                                                                 //      (terminated)
		.arqos                  (4'b0000),                                                                 //      (terminated)
		.awregion               (4'b0000),                                                                 //      (terminated)
		.arregion               (4'b0000),                                                                 //      (terminated)
		.wuser                  (8'b00000000),                                                             //      (terminated)
		.ruser                  (),                                                                        //      (terminated)
		.buser                  ()                                                                         //      (terminated)
	);

	altera_merlin_axi_translator #(
		.USE_S0_AWID                       (1),
		.USE_S0_AWREGION                   (0),
		.USE_M0_AWREGION                   (1),
		.USE_S0_AWLEN                      (1),
		.USE_S0_AWSIZE                     (1),
		.USE_S0_AWBURST                    (1),
		.USE_S0_AWLOCK                     (1),
		.USE_M0_AWLOCK                     (1),
		.USE_S0_AWCACHE                    (1),
		.USE_M0_AWCACHE                    (1),
		.USE_M0_AWPROT                     (1),
		.USE_S0_AWQOS                      (0),
		.USE_M0_AWQOS                      (1),
		.USE_S0_WSTRB                      (1),
		.USE_M0_WLAST                      (1),
		.USE_S0_BID                        (1),
		.USE_S0_BRESP                      (1),
		.USE_M0_BRESP                      (1),
		.USE_S0_ARID                       (1),
		.USE_S0_ARREGION                   (0),
		.USE_M0_ARREGION                   (1),
		.USE_S0_ARLEN                      (1),
		.USE_S0_ARSIZE                     (1),
		.USE_S0_ARBURST                    (1),
		.USE_S0_ARLOCK                     (1),
		.USE_M0_ARLOCK                     (1),
		.USE_M0_ARCACHE                    (1),
		.USE_M0_ARQOS                      (1),
		.USE_M0_ARPROT                     (1),
		.USE_S0_ARCACHE                    (1),
		.USE_S0_ARQOS                      (0),
		.USE_S0_RID                        (1),
		.USE_S0_RRESP                      (1),
		.USE_M0_RRESP                      (1),
		.USE_S0_RLAST                      (1),
		.M0_ID_WIDTH                       (2),
		.DATA_WIDTH                        (64),
		.S0_ID_WIDTH                       (12),
		.M0_ADDR_WIDTH                     (30),
		.S0_WRITE_ADDR_USER_WIDTH          (1),
		.S0_READ_ADDR_USER_WIDTH           (1),
		.M0_WRITE_ADDR_USER_WIDTH          (5),
		.M0_READ_ADDR_USER_WIDTH           (5),
		.S0_WRITE_DATA_USER_WIDTH          (1),
		.S0_WRITE_RESPONSE_DATA_USER_WIDTH (1),
		.S0_READ_DATA_USER_WIDTH           (1),
		.M0_WRITE_DATA_USER_WIDTH          (1),
		.M0_WRITE_RESPONSE_DATA_USER_WIDTH (1),
		.M0_READ_DATA_USER_WIDTH           (1),
		.S0_ADDR_WIDTH                     (30),
		.USE_S0_AWUSER                     (0),
		.USE_S0_ARUSER                     (0),
		.USE_S0_WUSER                      (0),
		.USE_S0_RUSER                      (0),
		.USE_S0_BUSER                      (0),
		.USE_M0_AWUSER                     (1),
		.USE_M0_ARUSER                     (1),
		.USE_M0_WUSER                      (0),
		.USE_M0_RUSER                      (0),
		.USE_M0_BUSER                      (0),
		.M0_AXI_VERSION                    ("AXI3"),
		.M0_BURST_LENGTH_WIDTH             (4),
		.S0_BURST_LENGTH_WIDTH             (4),
		.M0_LOCK_WIDTH                     (2),
		.S0_LOCK_WIDTH                     (2),
		.S0_AXI_VERSION                    ("AXI3")
	) id_pad (
		.aclk        (clk_clk),                                                              //       clk.clk
		.aresetn     (~rst_controller_reset_out_reset),                                      // clk_reset.reset_n
		.s0_awid     (hps_0_h2f_axi_master_awid),                                            //        s0.awid
		.s0_awaddr   (hps_0_h2f_axi_master_awaddr),                                          //          .awaddr
		.s0_awlen    (hps_0_h2f_axi_master_awlen),                                           //          .awlen
		.s0_awsize   (hps_0_h2f_axi_master_awsize),                                          //          .awsize
		.s0_awburst  (hps_0_h2f_axi_master_awburst),                                         //          .awburst
		.s0_awlock   (hps_0_h2f_axi_master_awlock),                                          //          .awlock
		.s0_awcache  (hps_0_h2f_axi_master_awcache),                                         //          .awcache
		.s0_awprot   (hps_0_h2f_axi_master_awprot),                                          //          .awprot
		.s0_awvalid  (hps_0_h2f_axi_master_awvalid),                                         //          .awvalid
		.s0_awready  (hps_0_h2f_axi_master_awready),                                         //          .awready
		.s0_wid      (hps_0_h2f_axi_master_wid),                                             //          .wid
		.s0_wdata    (hps_0_h2f_axi_master_wdata),                                           //          .wdata
		.s0_wstrb    (hps_0_h2f_axi_master_wstrb),                                           //          .wstrb
		.s0_wlast    (hps_0_h2f_axi_master_wlast),                                           //          .wlast
		.s0_wvalid   (hps_0_h2f_axi_master_wvalid),                                          //          .wvalid
		.s0_wready   (hps_0_h2f_axi_master_wready),                                          //          .wready
		.s0_bid      (hps_0_h2f_axi_master_bid),                                             //          .bid
		.s0_bresp    (hps_0_h2f_axi_master_bresp),                                           //          .bresp
		.s0_bvalid   (hps_0_h2f_axi_master_bvalid),                                          //          .bvalid
		.s0_bready   (hps_0_h2f_axi_master_bready),                                          //          .bready
		.s0_arid     (hps_0_h2f_axi_master_arid),                                            //          .arid
		.s0_araddr   (hps_0_h2f_axi_master_araddr),                                          //          .araddr
		.s0_arlen    (hps_0_h2f_axi_master_arlen),                                           //          .arlen
		.s0_arsize   (hps_0_h2f_axi_master_arsize),                                          //          .arsize
		.s0_arburst  (hps_0_h2f_axi_master_arburst),                                         //          .arburst
		.s0_arlock   (hps_0_h2f_axi_master_arlock),                                          //          .arlock
		.s0_arcache  (hps_0_h2f_axi_master_arcache),                                         //          .arcache
		.s0_arprot   (hps_0_h2f_axi_master_arprot),                                          //          .arprot
		.s0_arvalid  (hps_0_h2f_axi_master_arvalid),                                         //          .arvalid
		.s0_arready  (hps_0_h2f_axi_master_arready),                                         //          .arready
		.s0_rid      (hps_0_h2f_axi_master_rid),                                             //          .rid
		.s0_rdata    (hps_0_h2f_axi_master_rdata),                                           //          .rdata
		.s0_rresp    (hps_0_h2f_axi_master_rresp),                                           //          .rresp
		.s0_rlast    (hps_0_h2f_axi_master_rlast),                                           //          .rlast
		.s0_rvalid   (hps_0_h2f_axi_master_rvalid),                                          //          .rvalid
		.s0_rready   (hps_0_h2f_axi_master_rready),                                          //          .rready
		.m0_awid     (id_pad_m0_awid),                                                       //        m0.awid
		.m0_awaddr   (id_pad_m0_awaddr),                                                     //          .awaddr
		.m0_awlen    (id_pad_m0_awlen),                                                      //          .awlen
		.m0_awsize   (id_pad_m0_awsize),                                                     //          .awsize
		.m0_awburst  (id_pad_m0_awburst),                                                    //          .awburst
		.m0_awlock   (id_pad_m0_awlock),                                                     //          .awlock
		.m0_awcache  (id_pad_m0_awcache),                                                    //          .awcache
		.m0_awprot   (id_pad_m0_awprot),                                                     //          .awprot
		.m0_awuser   (id_pad_m0_awuser),                                                     //          .awuser
		.m0_awvalid  (id_pad_m0_awvalid),                                                    //          .awvalid
		.m0_awready  (id_pad_m0_awready),                                                    //          .awready
		.m0_wid      (id_pad_m0_wid),                                                        //          .wid
		.m0_wdata    (id_pad_m0_wdata),                                                      //          .wdata
		.m0_wstrb    (id_pad_m0_wstrb),                                                      //          .wstrb
		.m0_wlast    (id_pad_m0_wlast),                                                      //          .wlast
		.m0_wvalid   (id_pad_m0_wvalid),                                                     //          .wvalid
		.m0_wready   (id_pad_m0_wready),                                                     //          .wready
		.m0_bid      (id_pad_m0_bid),                                                        //          .bid
		.m0_bresp    (id_pad_m0_bresp),                                                      //          .bresp
		.m0_bvalid   (id_pad_m0_bvalid),                                                     //          .bvalid
		.m0_bready   (id_pad_m0_bready),                                                     //          .bready
		.m0_arid     (id_pad_m0_arid),                                                       //          .arid
		.m0_araddr   (id_pad_m0_araddr),                                                     //          .araddr
		.m0_arlen    (id_pad_m0_arlen),                                                      //          .arlen
		.m0_arsize   (id_pad_m0_arsize),                                                     //          .arsize
		.m0_arburst  (id_pad_m0_arburst),                                                    //          .arburst
		.m0_arlock   (id_pad_m0_arlock),                                                     //          .arlock
		.m0_arcache  (id_pad_m0_arcache),                                                    //          .arcache
		.m0_arprot   (id_pad_m0_arprot),                                                     //          .arprot
		.m0_aruser   (id_pad_m0_aruser),                                                     //          .aruser
		.m0_arvalid  (id_pad_m0_arvalid),                                                    //          .arvalid
		.m0_arready  (id_pad_m0_arready),                                                    //          .arready
		.m0_rid      (id_pad_m0_rid),                                                        //          .rid
		.m0_rdata    (id_pad_m0_rdata),                                                      //          .rdata
		.m0_rresp    (id_pad_m0_rresp),                                                      //          .rresp
		.m0_rlast    (id_pad_m0_rlast),                                                      //          .rlast
		.m0_rvalid   (id_pad_m0_rvalid),                                                     //          .rvalid
		.m0_rready   (id_pad_m0_rready),                                                     //          .rready
		.s0_awuser   (1'b0),                                                                 // (terminated)
		.s0_aruser   (1'b0),                                                                 // (terminated)
		.s0_awqos    (4'b0000),                                                              // (terminated)
		.s0_arqos    (4'b0000),                                                              // (terminated)
		.s0_awregion (4'b0000),                                                              // (terminated)
		.s0_arregion (4'b0000),                                                              // (terminated)
		.s0_wuser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_ruser    (),                                                                     // (terminated)
		.s0_buser    (),                                                                     // (terminated)
		.m0_awqos    (),                                                                     // (terminated)
		.m0_arqos    (),                                                                     // (terminated)
		.m0_awregion (),                                                                     // (terminated)
		.m0_arregion (),                                                                     // (terminated)
		.m0_wuser    (),                                                                     // (terminated)
		.m0_ruser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.m0_buser    (64'b0000000000000000000000000000000000000000000000000000000000000000)  // (terminated)
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (2),
		.ADDR_WIDTH                (30),
		.RDATA_WIDTH               (64),
		.WDATA_WIDTH               (64),
		.ADDR_USER_WIDTH           (5),
		.DATA_USER_WIDTH           (1),
		.AXI_BURST_LENGTH_WIDTH    (4),
		.AXI_LOCK_WIDTH            (2),
		.AXI_VERSION               ("AXI3"),
		.WRITE_ISSUING_CAPABILITY  (16),
		.READ_ISSUING_CAPABILITY   (16),
		.PKT_BEGIN_BURST           (135),
		.PKT_CACHE_H               (147),
		.PKT_CACHE_L               (144),
		.PKT_ADDR_SIDEBAND_H       (133),
		.PKT_ADDR_SIDEBAND_L       (129),
		.PKT_PROTECTION_H          (143),
		.PKT_PROTECTION_L          (141),
		.PKT_BURST_SIZE_H          (126),
		.PKT_BURST_SIZE_L          (124),
		.PKT_BURST_TYPE_H          (128),
		.PKT_BURST_TYPE_L          (127),
		.PKT_RESPONSE_STATUS_L     (148),
		.PKT_RESPONSE_STATUS_H     (149),
		.PKT_BURSTWRAP_H           (123),
		.PKT_BURSTWRAP_L           (116),
		.PKT_BYTE_CNT_H            (115),
		.PKT_BYTE_CNT_L            (108),
		.PKT_ADDR_H                (101),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_EXCLUSIVE       (107),
		.PKT_TRANS_LOCK            (106),
		.PKT_TRANS_COMPRESSED_READ (102),
		.PKT_TRANS_POSTED          (103),
		.PKT_TRANS_WRITE           (104),
		.PKT_TRANS_READ            (105),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (137),
		.PKT_SRC_ID_L              (137),
		.PKT_DEST_ID_H             (138),
		.PKT_DEST_ID_L             (138),
		.PKT_THREAD_ID_H           (140),
		.PKT_THREAD_ID_L           (139),
		.PKT_QOS_L                 (136),
		.PKT_QOS_H                 (136),
		.PKT_DATA_SIDEBAND_H       (134),
		.PKT_DATA_SIDEBAND_L       (134),
		.ST_DATA_W                 (150),
		.ST_CHANNEL_W              (2),
		.ID                        (0)
	) id_pad_m0_agent (
		.aclk                   (clk_clk),                                //              clk.clk
		.aresetn                (~rst_controller_reset_out_reset),        //        clk_reset.reset_n
		.write_cp_valid         (id_pad_m0_agent_write_cp_valid),         //         write_cp.valid
		.write_cp_data          (id_pad_m0_agent_write_cp_data),          //                 .data
		.write_cp_startofpacket (id_pad_m0_agent_write_cp_startofpacket), //                 .startofpacket
		.write_cp_endofpacket   (id_pad_m0_agent_write_cp_endofpacket),   //                 .endofpacket
		.write_cp_ready         (id_pad_m0_agent_write_cp_ready),         //                 .ready
		.write_rp_valid         (rsp_xbar_demux_src0_valid),              //         write_rp.valid
		.write_rp_data          (rsp_xbar_demux_src0_data),               //                 .data
		.write_rp_channel       (rsp_xbar_demux_src0_channel),            //                 .channel
		.write_rp_startofpacket (rsp_xbar_demux_src0_startofpacket),      //                 .startofpacket
		.write_rp_endofpacket   (rsp_xbar_demux_src0_endofpacket),        //                 .endofpacket
		.write_rp_ready         (rsp_xbar_demux_src0_ready),              //                 .ready
		.read_cp_valid          (id_pad_m0_agent_read_cp_valid),          //          read_cp.valid
		.read_cp_data           (id_pad_m0_agent_read_cp_data),           //                 .data
		.read_cp_startofpacket  (id_pad_m0_agent_read_cp_startofpacket),  //                 .startofpacket
		.read_cp_endofpacket    (id_pad_m0_agent_read_cp_endofpacket),    //                 .endofpacket
		.read_cp_ready          (id_pad_m0_agent_read_cp_ready),          //                 .ready
		.read_rp_valid          (rsp_xbar_demux_001_src0_valid),          //          read_rp.valid
		.read_rp_data           (rsp_xbar_demux_001_src0_data),           //                 .data
		.read_rp_channel        (rsp_xbar_demux_001_src0_channel),        //                 .channel
		.read_rp_startofpacket  (rsp_xbar_demux_001_src0_startofpacket),  //                 .startofpacket
		.read_rp_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),    //                 .endofpacket
		.read_rp_ready          (rsp_xbar_demux_001_src0_ready),          //                 .ready
		.awid                   (id_pad_m0_awid),                         // altera_axi_slave.awid
		.awaddr                 (id_pad_m0_awaddr),                       //                 .awaddr
		.awlen                  (id_pad_m0_awlen),                        //                 .awlen
		.awsize                 (id_pad_m0_awsize),                       //                 .awsize
		.awburst                (id_pad_m0_awburst),                      //                 .awburst
		.awlock                 (id_pad_m0_awlock),                       //                 .awlock
		.awcache                (id_pad_m0_awcache),                      //                 .awcache
		.awprot                 (id_pad_m0_awprot),                       //                 .awprot
		.awuser                 (id_pad_m0_awuser),                       //                 .awuser
		.awvalid                (id_pad_m0_awvalid),                      //                 .awvalid
		.awready                (id_pad_m0_awready),                      //                 .awready
		.wid                    (id_pad_m0_wid),                          //                 .wid
		.wdata                  (id_pad_m0_wdata),                        //                 .wdata
		.wstrb                  (id_pad_m0_wstrb),                        //                 .wstrb
		.wlast                  (id_pad_m0_wlast),                        //                 .wlast
		.wvalid                 (id_pad_m0_wvalid),                       //                 .wvalid
		.wready                 (id_pad_m0_wready),                       //                 .wready
		.bid                    (id_pad_m0_bid),                          //                 .bid
		.bresp                  (id_pad_m0_bresp),                        //                 .bresp
		.bvalid                 (id_pad_m0_bvalid),                       //                 .bvalid
		.bready                 (id_pad_m0_bready),                       //                 .bready
		.arid                   (id_pad_m0_arid),                         //                 .arid
		.araddr                 (id_pad_m0_araddr),                       //                 .araddr
		.arlen                  (id_pad_m0_arlen),                        //                 .arlen
		.arsize                 (id_pad_m0_arsize),                       //                 .arsize
		.arburst                (id_pad_m0_arburst),                      //                 .arburst
		.arlock                 (id_pad_m0_arlock),                       //                 .arlock
		.arcache                (id_pad_m0_arcache),                      //                 .arcache
		.arprot                 (id_pad_m0_arprot),                       //                 .arprot
		.aruser                 (id_pad_m0_aruser),                       //                 .aruser
		.arvalid                (id_pad_m0_arvalid),                      //                 .arvalid
		.arready                (id_pad_m0_arready),                      //                 .arready
		.rid                    (id_pad_m0_rid),                          //                 .rid
		.rdata                  (id_pad_m0_rdata),                        //                 .rdata
		.rresp                  (id_pad_m0_rresp),                        //                 .rresp
		.rlast                  (id_pad_m0_rlast),                        //                 .rlast
		.rvalid                 (id_pad_m0_rvalid),                       //                 .rvalid
		.rready                 (id_pad_m0_rready),                       //                 .rready
		.awqos                  (4'b0000),                                //      (terminated)
		.arqos                  (4'b0000),                                //      (terminated)
		.awregion               (4'b0000),                                //      (terminated)
		.arregion               (4'b0000),                                //      (terminated)
		.wuser                  (1'b0),                                   //      (terminated)
		.ruser                  (),                                       //      (terminated)
		.buser                  ()                                        //      (terminated)
	);

	altera_merlin_axi_slave_ni #(
		.PKT_QOS_H                   (100),
		.PKT_QOS_L                   (100),
		.PKT_THREAD_ID_H             (104),
		.PKT_THREAD_ID_L             (103),
		.PKT_RESPONSE_STATUS_H       (113),
		.PKT_RESPONSE_STATUS_L       (112),
		.PKT_BEGIN_BURST             (99),
		.PKT_CACHE_H                 (111),
		.PKT_CACHE_L                 (108),
		.PKT_DATA_SIDEBAND_H         (98),
		.PKT_DATA_SIDEBAND_L         (98),
		.PKT_ADDR_SIDEBAND_H         (97),
		.PKT_ADDR_SIDEBAND_L         (93),
		.PKT_BURST_TYPE_H            (92),
		.PKT_BURST_TYPE_L            (91),
		.PKT_PROTECTION_H            (107),
		.PKT_PROTECTION_L            (105),
		.PKT_BURST_SIZE_H            (90),
		.PKT_BURST_SIZE_L            (88),
		.PKT_BURSTWRAP_H             (87),
		.PKT_BURSTWRAP_L             (80),
		.PKT_BYTE_CNT_H              (79),
		.PKT_BYTE_CNT_L              (72),
		.PKT_ADDR_H                  (65),
		.PKT_ADDR_L                  (36),
		.PKT_TRANS_EXCLUSIVE         (71),
		.PKT_TRANS_LOCK              (70),
		.PKT_TRANS_COMPRESSED_READ   (66),
		.PKT_TRANS_POSTED            (67),
		.PKT_TRANS_WRITE             (68),
		.PKT_TRANS_READ              (69),
		.PKT_DATA_H                  (31),
		.PKT_DATA_L                  (0),
		.PKT_BYTEEN_H                (35),
		.PKT_BYTEEN_L                (32),
		.PKT_SRC_ID_H                (101),
		.PKT_SRC_ID_L                (101),
		.PKT_DEST_ID_H               (102),
		.PKT_DEST_ID_L               (102),
		.ADDR_USER_WIDTH             (5),
		.DATA_USER_WIDTH             (1),
		.ST_DATA_W                   (114),
		.ADDR_WIDTH                  (30),
		.RDATA_WIDTH                 (32),
		.WDATA_WIDTH                 (32),
		.ST_CHANNEL_W                (2),
		.AXI_SLAVE_ID_W              (2),
		.PASS_ID_TO_SLAVE            (1),
		.AXI_VERSION                 ("AXI3"),
		.WRITE_ACCEPTANCE_CAPABILITY (1),
		.READ_ACCEPTANCE_CAPABILITY  (1)
	) merlin_axi_master_ni_0_altera_axi_slave_agent (
		.aclk                   (clk_clk),                                                                 //        clock_sink.clk
		.aresetn                (~rst_controller_reset_out_reset),                                         //        reset_sink.reset_n
		.read_cp_valid          (burst_adapter_001_source0_valid),                                         //           read_cp.valid
		.read_cp_ready          (burst_adapter_001_source0_ready),                                         //                  .ready
		.read_cp_data           (burst_adapter_001_source0_data),                                          //                  .data
		.read_cp_channel        (burst_adapter_001_source0_channel),                                       //                  .channel
		.read_cp_startofpacket  (burst_adapter_001_source0_startofpacket),                                 //                  .startofpacket
		.read_cp_endofpacket    (burst_adapter_001_source0_endofpacket),                                   //                  .endofpacket
		.write_cp_ready         (burst_adapter_source0_ready),                                             //          write_cp.ready
		.write_cp_valid         (burst_adapter_source0_valid),                                             //                  .valid
		.write_cp_data          (burst_adapter_source0_data),                                              //                  .data
		.write_cp_channel       (burst_adapter_source0_channel),                                           //                  .channel
		.write_cp_startofpacket (burst_adapter_source0_startofpacket),                                     //                  .startofpacket
		.write_cp_endofpacket   (burst_adapter_source0_endofpacket),                                       //                  .endofpacket
		.read_rp_ready          (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_ready),             //           read_rp.ready
		.read_rp_valid          (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_valid),             //                  .valid
		.read_rp_data           (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_data),              //                  .data
		.read_rp_startofpacket  (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_startofpacket),     //                  .startofpacket
		.read_rp_endofpacket    (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_endofpacket),       //                  .endofpacket
		.write_rp_ready         (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_ready),            //          write_rp.ready
		.write_rp_valid         (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_valid),            //                  .valid
		.write_rp_data          (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_data),             //                  .data
		.write_rp_startofpacket (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_startofpacket),    //                  .startofpacket
		.write_rp_endofpacket   (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_endofpacket),      //                  .endofpacket
		.awid                   (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awid),    // altera_axi_master.awid
		.awaddr                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awaddr),  //                  .awaddr
		.awlen                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlen),   //                  .awlen
		.awsize                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awsize),  //                  .awsize
		.awburst                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awburst), //                  .awburst
		.awlock                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awlock),  //                  .awlock
		.awcache                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awcache), //                  .awcache
		.awprot                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awprot),  //                  .awprot
		.awuser                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awuser),  //                  .awuser
		.awvalid                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awvalid), //                  .awvalid
		.awready                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_awready), //                  .awready
		.wid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wid),     //                  .wid
		.wdata                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wdata),   //                  .wdata
		.wstrb                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wstrb),   //                  .wstrb
		.wlast                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wlast),   //                  .wlast
		.wvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wvalid),  //                  .wvalid
		.wready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_wready),  //                  .wready
		.bid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bid),     //                  .bid
		.bresp                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bresp),   //                  .bresp
		.bvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bvalid),  //                  .bvalid
		.bready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_bready),  //                  .bready
		.arid                   (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arid),    //                  .arid
		.araddr                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_araddr),  //                  .araddr
		.arlen                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlen),   //                  .arlen
		.arsize                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arsize),  //                  .arsize
		.arburst                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arburst), //                  .arburst
		.arlock                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arlock),  //                  .arlock
		.arcache                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arcache), //                  .arcache
		.arprot                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arprot),  //                  .arprot
		.aruser                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_aruser),  //                  .aruser
		.arvalid                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arvalid), //                  .arvalid
		.arready                (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_arready), //                  .arready
		.rid                    (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rid),     //                  .rid
		.rdata                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rdata),   //                  .rdata
		.rresp                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rresp),   //                  .rresp
		.rlast                  (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rlast),   //                  .rlast
		.rvalid                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rvalid),  //                  .rvalid
		.rready                 (merlin_axi_master_ni_0_altera_axi_slave_agent_altera_axi_master_rready)   //                  .rready
	);

	axi_agent_addr_router addr_router (
		.sink_ready         (id_pad_m0_agent_write_cp_ready),         //      sink.ready
		.sink_valid         (id_pad_m0_agent_write_cp_valid),         //          .valid
		.sink_data          (id_pad_m0_agent_write_cp_data),          //          .data
		.sink_startofpacket (id_pad_m0_agent_write_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (id_pad_m0_agent_write_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready          (addr_router_src_ready),                  //       src.ready
		.src_valid          (addr_router_src_valid),                  //          .valid
		.src_data           (addr_router_src_data),                   //          .data
		.src_channel        (addr_router_src_channel),                //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)             //          .endofpacket
	);

	axi_agent_addr_router addr_router_001 (
		.sink_ready         (id_pad_m0_agent_read_cp_ready),         //      sink.ready
		.sink_valid         (id_pad_m0_agent_read_cp_valid),         //          .valid
		.sink_data          (id_pad_m0_agent_read_cp_data),          //          .data
		.sink_startofpacket (id_pad_m0_agent_read_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (id_pad_m0_agent_read_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),             //       src.ready
		.src_valid          (addr_router_001_src_valid),             //          .valid
		.src_data           (addr_router_001_src_data),              //          .data
		.src_channel        (addr_router_001_src_channel),           //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),     //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)        //          .endofpacket
	);

	axi_agent_id_router id_router (
		.sink_ready         (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_ready),         //      sink.ready
		.sink_valid         (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_valid),         //          .valid
		.sink_data          (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_data),          //          .data
		.sink_startofpacket (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (merlin_axi_master_ni_0_altera_axi_slave_agent_write_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                  //          .valid
		.src_data           (id_router_src_data),                                                   //          .data
		.src_channel        (id_router_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                             //          .endofpacket
	);

	axi_agent_id_router id_router_001 (
		.sink_ready         (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_ready),         //      sink.ready
		.sink_valid         (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_valid),         //          .valid
		.sink_data          (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_data),          //          .data
		.sink_startofpacket (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (merlin_axi_master_ni_0_altera_axi_slave_agent_read_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                             //          .valid
		.src_data           (id_router_001_src_data),                                              //          .data
		.src_channel        (id_router_001_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (99),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (72),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (90),
		.PKT_BURST_SIZE_L          (88),
		.PKT_BURST_TYPE_H          (92),
		.PKT_BURST_TYPE_L          (91),
		.PKT_BURSTWRAP_H           (87),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.OUT_NARROW_SIZE           (1),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (1),
		.OUT_COMPLETE_WRAP         (1),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (78),
		.OUT_BURSTWRAP_H           (87),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter (
		.clk                   (clk_clk),                                //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),         // cr0_reset.reset
		.sink0_valid           (width_adapter_cmd_source_valid),         //     sink0.valid
		.sink0_data            (width_adapter_cmd_source_data),          //          .data
		.sink0_channel         (width_adapter_cmd_source_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_cmd_source_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_cmd_source_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_cmd_source_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),            //   source0.valid
		.source0_data          (burst_adapter_source0_data),             //          .data
		.source0_channel       (burst_adapter_source0_channel),          //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket),    //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),      //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)             //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (99),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (72),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (90),
		.PKT_BURST_SIZE_L          (88),
		.PKT_BURST_TYPE_H          (92),
		.PKT_BURST_TYPE_L          (91),
		.PKT_BURSTWRAP_H           (87),
		.PKT_BURSTWRAP_L           (80),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.OUT_NARROW_SIZE           (1),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (1),
		.OUT_COMPLETE_WRAP         (1),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (78),
		.OUT_BURSTWRAP_H           (87),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),             // cr0_reset.reset
		.sink0_valid           (width_adapter_001_cmd_source_valid),         //     sink0.valid
		.sink0_data            (width_adapter_001_cmd_source_data),          //          .data
		.sink0_channel         (width_adapter_001_cmd_source_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_001_cmd_source_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_001_cmd_source_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_001_cmd_source_ready),         //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),            //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),             //          .data
		.source0_channel       (burst_adapter_001_source0_channel),          //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket),    //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),      //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)             //          .ready
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (101),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (115),
		.IN_PKT_BYTE_CNT_L             (108),
		.IN_PKT_TRANS_COMPRESSED_READ  (102),
		.IN_PKT_BURSTWRAP_H            (123),
		.IN_PKT_BURSTWRAP_L            (116),
		.IN_PKT_BURST_SIZE_H           (126),
		.IN_PKT_BURST_SIZE_L           (124),
		.IN_PKT_RESPONSE_STATUS_H      (149),
		.IN_PKT_RESPONSE_STATUS_L      (148),
		.IN_PKT_TRANS_EXCLUSIVE        (107),
		.IN_PKT_BURST_TYPE_H           (128),
		.IN_PKT_BURST_TYPE_L           (127),
		.IN_PKT_TRANS_POSTED           (103),
		.IN_ST_DATA_W                  (150),
		.OUT_PKT_ADDR_H                (65),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (72),
		.OUT_PKT_TRANS_COMPRESSED_READ (66),
		.OUT_PKT_TRANS_EXCLUSIVE       (71),
		.OUT_PKT_RESPONSE_STATUS_H     (113),
		.OUT_PKT_RESPONSE_STATUS_L     (112),
		.OUT_PKT_BURST_SIZE_H          (90),
		.OUT_PKT_BURST_SIZE_L          (88),
		.OUT_PKT_BURST_TYPE_H          (92),
		.OUT_PKT_BURST_TYPE_L          (91),
		.OUT_ST_DATA_W                 (114),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter (
		.clk                   (clk_clk),                                //      clock.clk
		.reset                 (rst_controller_reset_out_reset),         //      reset.reset
		.cmd_in_valid          (cmd_xbar_demux_src0_valid),              //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_demux_src0_channel),            //           .channel
		.cmd_in_data           (cmd_xbar_demux_src0_data),               //           .data
		.cmd_in_startofpacket  (cmd_xbar_demux_src0_startofpacket),      //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_demux_src0_endofpacket),        //           .endofpacket
		.cmd_in_ready          (cmd_xbar_demux_src0_ready),              //           .ready
		.cmd_out_ready         (width_adapter_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_src_channel),                  //           .channel
		.rsp_in_data           (id_router_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (101),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (115),
		.IN_PKT_BYTE_CNT_L             (108),
		.IN_PKT_TRANS_COMPRESSED_READ  (102),
		.IN_PKT_BURSTWRAP_H            (123),
		.IN_PKT_BURSTWRAP_L            (116),
		.IN_PKT_BURST_SIZE_H           (126),
		.IN_PKT_BURST_SIZE_L           (124),
		.IN_PKT_RESPONSE_STATUS_H      (149),
		.IN_PKT_RESPONSE_STATUS_L      (148),
		.IN_PKT_TRANS_EXCLUSIVE        (107),
		.IN_PKT_BURST_TYPE_H           (128),
		.IN_PKT_BURST_TYPE_L           (127),
		.IN_PKT_TRANS_POSTED           (103),
		.IN_ST_DATA_W                  (150),
		.OUT_PKT_ADDR_H                (65),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (72),
		.OUT_PKT_TRANS_COMPRESSED_READ (66),
		.OUT_PKT_TRANS_EXCLUSIVE       (71),
		.OUT_PKT_RESPONSE_STATUS_H     (113),
		.OUT_PKT_RESPONSE_STATUS_L     (112),
		.OUT_PKT_BURST_SIZE_H          (90),
		.OUT_PKT_BURST_SIZE_L          (88),
		.OUT_PKT_BURST_TYPE_H          (92),
		.OUT_PKT_BURST_TYPE_L          (91),
		.OUT_ST_DATA_W                 (114),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter_001 (
		.clk                   (clk_clk),                                    //      clock.clk
		.reset                 (rst_controller_reset_out_reset),             //      reset.reset
		.cmd_in_valid          (cmd_xbar_demux_001_src0_valid),              //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_demux_001_src0_channel),            //           .channel
		.cmd_in_data           (cmd_xbar_demux_001_src0_data),               //           .data
		.cmd_in_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),      //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),        //           .endofpacket
		.cmd_in_ready          (cmd_xbar_demux_001_src0_ready),              //           .ready
		.cmd_out_ready         (width_adapter_001_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_001_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_001_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_001_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_001_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_001_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_001_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_001_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_001_src_channel),                  //           .channel
		.rsp_in_data           (id_router_001_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_001_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_001_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_001_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_001_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_001_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_001_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_001_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_001_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	axi_agent_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	axi_agent_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	axi_agent_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready         (width_adapter_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)         //          .endofpacket
	);

	axi_agent_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),             // clk_reset.reset
		.sink_ready         (width_adapter_001_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_001_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_001_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)         //          .endofpacket
	);

endmodule
